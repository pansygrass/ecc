`timescale 1 ns /1 ps

module dec_tb();

reg [74:0] IN;
wire [62:0] OUT;
wire [11:0] SYN;
wire ERR, SGL, DBL;
reg clk;

// Fake clock does nothing
dec_top DUT0 (.IN(IN), .OUT(OUT), .SYN(SYN), .ERR(ERR), .SGL(SGL), .DBL(DBL), .clk(clk));
initial begin

$vcdpluson;
    IN <= 75'd0;
    #`CLOCK_PERIOD IN <= 75'b000000000000000000000000000000000000000000000000000000000000000000000000000; 
    #`CLOCK_PERIOD IN <= 75'b010100111001000000000000000000000000000000000000000000000000000000000000001;
    #`CLOCK_PERIOD IN <= 75'b010100111001000000000000000000000000000000000000000000000000000000000000011;
    #`CLOCK_PERIOD IN <= 75'b010100111001000000000000000000000000000000000000000000000000000000000000111;
    #`CLOCK_PERIOD IN <= 75'b010100111001000000000000000000000000000000000000000000000000000000000001111;
    #`CLOCK_PERIOD IN <= 75'b101001110010000000000000000000000000000000000000000000000000000000000000010;
    #`CLOCK_PERIOD IN <= 75'b111101001011000000000000000000000000000000000000000000000000000000000000011;
    #`CLOCK_PERIOD IN <= 75'b000111011101000000000000000000000000000000000000000000000000000000000000100;
    #`CLOCK_PERIOD IN <= 75'b010011100100000000000000000000000000000000000000000000000000000000000000101;
    #`CLOCK_PERIOD IN <= 75'b101110101111000000000000000000000000000000000000000000000000000000000000110;
    #`CLOCK_PERIOD IN <= 75'b111010010110000000000000000000000000000000000000000000000000000000000000111;
    #`CLOCK_PERIOD IN <= 75'b001110111010000000000000000000000000000000000000000000000000000000000001000;
    #`CLOCK_PERIOD IN <= 75'b011010000011000000000000000000000000000000000000000000000000000000000001001;
$vcdplusoff;

end

initial begin
    $monitor($time, ": IN=%b, OUT=%b, SYN=%b, ERR=%b, SGL=%b, DBL=%b", IN, OUT, SYN, ERR, SGL, DBL);
end

endmodule

