`timescale 1 ns /1 ps

module dec_tb();

reg [140:0] IN;
wire [126:0] OUT;
wire [13:0] SYN;
wire ERR, SGL, DBL;
reg clk;

// Fake clock does nothing
dec_top DUT0 (.IN(IN), .OUT(OUT), .SYN(SYN), .ERR(ERR), .SGL(SGL), .DBL(DBL), .clk(clk));
initial begin

$vcdpluson;
    IN <= 141'd0;
    #`CLOCK_PERIOD IN <= 141'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    #`CLOCK_PERIOD IN <= 141'b000011011101110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001;
    #`CLOCK_PERIOD IN <= 141'b000011011101110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011;
    #`CLOCK_PERIOD IN <= 141'b000011011101110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111;
    #`CLOCK_PERIOD IN <= 141'b000011011101110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111;
    #`CLOCK_PERIOD IN <= 141'b000110111011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010;
    #`CLOCK_PERIOD IN <= 141'b000101100110010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011;
    #`CLOCK_PERIOD IN <= 141'b001101110111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100;
    #`CLOCK_PERIOD IN <= 141'b001110101010110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101;
    #`CLOCK_PERIOD IN <= 141'b001011001100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110;
    #`CLOCK_PERIOD IN <= 141'b001000010001010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111;
    #`CLOCK_PERIOD IN <= 141'b011011101110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000;
    #`CLOCK_PERIOD IN <= 141'b011000110011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001;
$vcdplusoff;

end

initial begin
    $monitor($time, ": IN=%b, OUT=%b, SYN=%b, ERR=%b, SGL=%b, DBL=%b", IN, OUT, SYN, ERR, SGL, DBL);
end

endmodule

