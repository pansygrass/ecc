`timescale 1 ns /1 ps

module dec_tb();

reg [40:0] IN;
wire [30:0] OUT;
wire [9:0] SYN;
wire ERR, SGL, DBL;
reg clk;

// Fake clock does nothing
dec_top DUT0 (.IN(IN), .OUT(OUT), .SYN(SYN), .ERR(ERR), .SGL(SGL), .DBL(DBL), .clk(clk));
initial begin
$vcdpluson;
    IN <= 41'd0;
    #`CLOCK_PERIOD IN <= 41'b00000000000000000000000000000000000000000; 
    #`CLOCK_PERIOD IN <= 41'b11110001101110101111110110011101001111000;
    #`CLOCK_PERIOD IN <= 41'b11101000100111100001101101101010000010101;
    #`CLOCK_PERIOD IN <= 41'b00010011001010110011011110000111001010110;
    #`CLOCK_PERIOD IN <= 41'b10000101111100010110101111110011001101100;
    #`CLOCK_PERIOD IN <= 41'b00011101101001111100011101011000101000101;
    #`CLOCK_PERIOD IN <= 41'b01010011111111110100001101000110100001101;
    #`CLOCK_PERIOD IN <= 41'b00110011000101010001011110010001010010000;
    #`CLOCK_PERIOD IN <= 41'b01000000100010110010011101111111011000101;
    #`CLOCK_PERIOD IN <= 41'b00111110100000011011001001111011010011110;
    #`CLOCK_PERIOD IN <= 41'b10011001011010101001110110110010011100101;
$vcdplusoff;

end

initial begin
    $monitor($time, ": IN=%b, OUT=%b, SYN=%b, ERR=%b, SGL=%b, DBL=%b", IN, OUT, SYN, ERR, SGL, DBL);
end

endmodule


