`timescale 1 ns /1 ps

module dec_tb();

reg [71:0] IN;
wire [71:0] OUT;
wire [7:0] SYN;
wire ERR, SGL, DBL;
reg clk;

// Fake clock does nothing
dec_top DUT0 (.IN(IN), .OUT(OUT), .SYN(SYN), .ERR(ERR), .SGL(SGL), .DBL(DBL), .clk(clk));
initial begin

$vcdpluson;
    IN <= 72'd0;
    #`CLOCK_PERIOD IN <= 72'b000000000000000000000000000000000000000000000000000000000000000000000000;
    #`CLOCK_PERIOD IN <= 72'b000000000000000000000010000000100000000000000000000000000000000000000000;
    #`CLOCK_PERIOD IN <= 72'b001000110000000000000000000000000000000000000000000000000000000000000001;
    #`CLOCK_PERIOD IN <= 72'b001010110000000000000000000000000000000000000000000000000000000000000001;
    #`CLOCK_PERIOD IN <= 72'b010000110000000000000000000000000000000000000000000000000000000000000010;
    #`CLOCK_PERIOD IN <= 72'b011000000000000000000000000000000000000000000000000000000000000000000011;
    #`CLOCK_PERIOD IN <= 72'b100000110000000000000000000000000000000000000000000000000000000000000100;
    #`CLOCK_PERIOD IN <= 72'b101000000000000000000000000000000000000000000000000000000000000000000101;
    #`CLOCK_PERIOD IN <= 72'b110000000000000000000000000000000000000000000000000000000000000000000110;
    #`CLOCK_PERIOD IN <= 72'b111000110000000000000000000000000000000000000000000000000000000000000111;
    #`CLOCK_PERIOD IN <= 72'b001111010000000000000000000000000000000000000000000000000000000000001000;
    #`CLOCK_PERIOD IN <= 72'b000111100000000000000000000000000000000000000000000000000000000000001001;
$vcdplusoff;

end

initial begin
    $monitor($time, ": IN=%b, OUT=%b, SYN=%b, ERR=%b, SGL=%b, DBL=%b", IN, OUT, SYN, ERR, SGL, DBL);
end

endmodule

