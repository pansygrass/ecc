`timescale 1 ns /1 ps

module dec_tb();

reg [71:0] IN;
wire [71:0] OUT;
wire [7:0] SYN;
wire ERR, SGL, DBL;
reg clk;

// Fake clock does nothing
dec_top DUT0 (.IN(IN), .OUT(OUT), .SYN(SYN), .ERR(ERR), .SGL(SGL), .DBL(DBL), .clk(clk));
initial begin

$vcdpluson;
    IN <= 72'd0;
    #`CLOCK_PERIOD IN <= 72'b000000000000000000000000000000000000000000000000000000000000000000000000;
    #`CLOCK_PERIOD IN <= 72'b010110100001000111000110110000110101000100001101110000001000001000011000;
    #`CLOCK_PERIOD IN <= 72'b001001100010110110111011001100000110111100010000111001011111001110111111;
    #`CLOCK_PERIOD IN <= 72'b101100110110010000100110000100101011010000010111010000000011110010110001;
    #`CLOCK_PERIOD IN <= 72'b101111000100111001011100111110011111100111100000100000011000001110000101;
    #`CLOCK_PERIOD IN <= 72'b000011110100001100011001101111001010001001001111000000000101011010011101;
    #`CLOCK_PERIOD IN <= 72'b111100110101011111100011110111000000111001111001010011100000001000101110;
    #`CLOCK_PERIOD IN <= 72'b100100010110101010101001110100001101010010100000110001011100111001011101;
    #`CLOCK_PERIOD IN <= 72'b000001100011100000111010101111011011000100111001011101001111101111101011;
    #`CLOCK_PERIOD IN <= 72'b111001110110110100000100111110010000100110011101110110001100100000011000;
$vcdplusoff;

end

initial begin
    $monitor($time, ": IN=%b, OUT=%b, SYN=%b, ERR=%b, SGL=%b, DBL=%b", IN, OUT, SYN, ERR, SGL, DBL);
end

endmodule

