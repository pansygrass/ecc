`timescale 1 ns /1 ps

module dec_tb();

reg [74:0] IN;
wire [62:0] OUT;
wire [11:0] SYN;
wire ERR, SGL, DBL;
reg clk;

// Fake clock does nothing
dec_top DUT0 (.IN(IN), .OUT(OUT), .SYN(SYN), .ERR(ERR), .SGL(SGL), .DBL(DBL), .clk(clk));
initial begin

$vcdpluson;
    IN <= 75'd0;
    #`CLOCK_PERIOD IN <= 75'b000000000000000000000000000000000000000000000000000000000000000000000000000; 
    #`CLOCK_PERIOD IN <= 75'b101111110001001000111000110110000110101000100001101110000001000001000011000;
    #`CLOCK_PERIOD IN <= 75'b111110110010010110110111011001100000110111100010000111001011111001110111111;
    #`CLOCK_PERIOD IN <= 75'b010111101000110010000100110000100101011010000010111010000000011110010110001;
    #`CLOCK_PERIOD IN <= 75'b001101001100100111001011100111110011111100111100000100000011000001110000101;
    #`CLOCK_PERIOD IN <= 75'b010000000110100001100011001101111001010001001001111000000000101011010011101;
    #`CLOCK_PERIOD IN <= 75'b101100011100101011111100011110111000000111001111001010011100000001000101110;
    #`CLOCK_PERIOD IN <= 75'b001101111011110101010101001110100001101010010100000110001011100111001011101;
    #`CLOCK_PERIOD IN <= 75'b111110101000011100000111010101111011011000100111001011101001111101111101011;
    #`CLOCK_PERIOD IN <= 75'b001000101001110110100000100111110010000100110011101110110001100100000011000;
$vcdplusoff;

end

initial begin
    $monitor($time, ": IN=%b, OUT=%b, SYN=%b, ERR=%b, SGL=%b, DBL=%b", IN, OUT, SYN, ERR, SGL, DBL);
end

endmodule

