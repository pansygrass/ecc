`timescale 1 ns /1 ps

module dec_tb();

reg [136:0] IN;
wire [136:0] OUT;
wire [8:0] SYN;
wire ERR, SGL, DBL;
reg clk;

// Fake clock does nothing
dec_top DUT0 (.IN(IN), .OUT(OUT), .SYN(SYN), .ERR(ERR), .SGL(SGL), .DBL(DBL), .clk(clk));
initial begin

$vcdpluson;
    IN <= 137'd0;

    #`CLOCK_PERIOD IN <= 137'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    #`CLOCK_PERIOD IN <= 137'b11100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001;
    #`CLOCK_PERIOD IN <= 137'b11100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011;
    #`CLOCK_PERIOD IN <= 137'b11100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111;
    #`CLOCK_PERIOD IN <= 137'b11010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010;
    #`CLOCK_PERIOD IN <= 137'b00110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011;
    #`CLOCK_PERIOD IN <= 137'b01110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100;
    #`CLOCK_PERIOD IN <= 137'b10010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101;
    #`CLOCK_PERIOD IN <= 137'b10100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110;
    #`CLOCK_PERIOD IN <= 137'b01000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111;
    #`CLOCK_PERIOD IN <= 137'b10110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000;
    #`CLOCK_PERIOD IN <= 137'b01010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001;
$vcdplusoff;

end

initial begin
    $monitor($time, ": IN=%b, OUT=%b, SYN=%b, ERR=%b, SGL=%b, DBL=%b", IN, OUT, SYN, ERR, SGL, DBL);
end

endmodule

