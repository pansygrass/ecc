`timescale 1 ns /1 ps

module dec_tb();

reg [140:0] IN;
wire [126:0] OUT;
wire [13:0] SYN;
wire ERR, SGL, DBL;
reg clk;

// Fake clock does nothing
dec_top DUT0 (.IN(IN), .OUT(OUT), .SYN(SYN), .ERR(ERR), .SGL(SGL), .DBL(DBL), .clk(clk));
initial begin

$vcdpluson;
    IN <= 141'd0;
    #`CLOCK_PERIOD IN <= 141'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    #`CLOCK_PERIOD IN <= 141'b010010001001001010011101101111110110000111111000101000000010001001010111100100010001001100010100110111000011100100010000110001010010100111111;
    #`CLOCK_PERIOD IN <= 141'b101111110111010000001110001001011110001000000110011111100010011101000101101100100010110011010001100110001111000000011011101001001011000110011;
    #`CLOCK_PERIOD IN <= 141'b110000001001100010111111011001100011110100000110101110011010000010101100111111000011000100110001100011000110100010000110011101110111111010001;
    #`CLOCK_PERIOD IN <= 141'b010001111111011010000100101001011011011000000111110110101011001111100000101001001011100100011101101101110101001101011100100110011100011010111;
    #`CLOCK_PERIOD IN <= 141'b001001011001011110000101011111010101011010010010001011011011011000110011011101111010101101111011100010010100110001101100000001001001011001010;
    #`CLOCK_PERIOD IN <= 141'b100101111101001100111010011001100011011100010110101010001011001110000111011011110110011010111101101011110110111110001001000000000001011110000;
    #`CLOCK_PERIOD IN <= 141'b001001010100110110101011011000100101010011101000101100100011000011001000110100100100010100110011111101011101011010011110010100011111000111000;
    #`CLOCK_PERIOD IN <= 141'b100001111010000010110100011111101110010111001001011001100010000010110000110111011001101000100001110101011011001110000011000110100100001110010;
    #`CLOCK_PERIOD IN <= 141'b000100111110111101000101000001011110010111010011100110111000011100110000010000110001101111111000000000100100001010101110011110111110110001111;
    #`CLOCK_PERIOD IN <= 141'b111010110001101010010110110011010101100001101001001101010011001000011101001101100011010011011111101111011110101001100110000100011110111111000;
$vcdplusoff;

end

initial begin
    $monitor($time, ": IN=%b, OUT=%b, SYN=%b, ERR=%b, SGL=%b, DBL=%b", IN, OUT, SYN, ERR, SGL, DBL);
end

endmodule

