`timescale 1 ns /1 ps

module dec_tb();

reg [38:0] IN;
wire [38:0] OUT;
wire [6:0] SYN;
wire ERR, SGL, DBL;
reg clk;

// Fake clock does nothing
dec_top DUT0 (.IN(IN), .OUT(OUT), .SYN(SYN), .ERR(ERR), .SGL(SGL), .DBL(DBL), .clk(clk));
initial begin

$vcdpluson;
    IN <= 32'd0;
    #`CLOCK_PERIOD IN <= 39'b000000000000000000000000000000000000011;
    #`CLOCK_PERIOD IN <= 39'b001111001110101111110110011101001111011;
    #`CLOCK_PERIOD IN <= 39'b001001100111100001101101101010000010110;
    #`CLOCK_PERIOD IN <= 39'b101101011010110011011110000111001010101;
    #`CLOCK_PERIOD IN <= 39'b011001101100010110101111110011001101111;
    #`CLOCK_PERIOD IN <= 39'b100101011001111100011101011000101000110;
    #`CLOCK_PERIOD IN <= 39'b001011011111110100001101000110100001110;
    #`CLOCK_PERIOD IN <= 39'b100011010101010001011110010001010010011;
    #`CLOCK_PERIOD IN <= 39'b000001100010110010011101111111011000110;
    #`CLOCK_PERIOD IN <= 39'b110110000000011011001001111011010011101;
    #`CLOCK_PERIOD IN <= 39'b010110001010101001110110110010011100110;
$vcdplusoff;

end

initial begin
    $monitor($time, ": IN=%b, OUT=%b, SYN=%b, ERR=%b, SGL=%b, DBL=%b", IN, OUT, SYN, ERR, SGL, DBL);
end

endmodule


//Original data, no errors
//000000000000000000000000000000000000000;
//001111001110101111110110011101001111000;
//001001100111100001101101101010000010101;
//101101011010110011011110000111001010110;
//011001101100010110101111110011001101100;
//100101011001111100011101011000101000101;
//001011011111110100001101000110100001101;
//100011010101010001011110010001010010000;
//000001100010110010011101111111011000101;
//110110000000011011001001111011010011110;
//010110001010101001110110110010011100101;
