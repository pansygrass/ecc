`timescale 1 ns /1 ps

module enc_top_tb();

reg [126:0] IN;
wire [140:0] OUT;
reg clk;

// Fake clock does nothing
enc_top DUT0 (.IN(IN), .OUT(OUT), .clk(clk));

initial begin

$vcdpluson;
    IN <= 127'd0;
    #`CLOCK_PERIOD IN <= 128'd111280905621495480921325258608442123583;
    #`CLOCK_PERIOD IN <= 128'd2350736407967074960062813466992612915  ;
    #`CLOCK_PERIOD IN <= 128'd31801674904286656728433206597602176977 ;
    #`CLOCK_PERIOD IN <= 128'd107110406285996782703011031750322370775;
    #`CLOCK_PERIOD IN <= 128'd149785652147276348631935800520558547658;
    #`CLOCK_PERIOD IN <= 128'd137309132015708669817313440322734260976;
    #`CLOCK_PERIOD IN <= 128'd71011365181347901178350486250909744696 ;
    #`CLOCK_PERIOD IN <= 128'd29989991159215892356985217153094600818 ;
    #`CLOCK_PERIOD IN <= 128'd139074306924167799490053291585714486671;
    #`CLOCK_PERIOD IN <= 128'd110126893406634927828874494532336631288;
$vcdplusoff;

end

initial begin
    $monitor($time, ": IN=%b, OUT=%b", IN, OUT);
end

endmodule

