`timescale 1 ns /1 ps

module dec_tb();

reg [40:0] IN;
wire [30:0] OUT;
wire [9:0] SYN;
wire ERR, SGL, DBL;
reg clk;

// Fake clock does nothing
dec_top DUT0 (.IN(IN), .OUT(OUT), .SYN(SYN), .ERR(ERR), .SGL(SGL), .DBL(DBL), .clk(clk));
initial begin
$vcdpluson;
    IN <= 41'd0;
    #`CLOCK_PERIOD IN <= 41'b00000000000000000000000000000000000000000; 
    #`CLOCK_PERIOD IN <= 41'b11011010010000000000000000000000000000001;
    #`CLOCK_PERIOD IN <= 41'b11011010010000000000000000000000000000011;
    #`CLOCK_PERIOD IN <= 41'b11011010010000000000000000000000000000111;
    #`CLOCK_PERIOD IN <= 41'b11011010010000000000000000000000000001111;
    #`CLOCK_PERIOD IN <= 41'b01101110110000000000000000000000000000010;
    #`CLOCK_PERIOD IN <= 41'b10110100100000000000000000000000000000011;
    #`CLOCK_PERIOD IN <= 41'b11011101100000000000000000000000000000100;
    #`CLOCK_PERIOD IN <= 41'b00000111110000000000000000000000000000101;
    #`CLOCK_PERIOD IN <= 41'b10110011010000000000000000000000000000110;
    #`CLOCK_PERIOD IN <= 41'b01101001000000000000000000000000000000111;
    #`CLOCK_PERIOD IN <= 41'b01100001010000000000000000000000000001000;
    #`CLOCK_PERIOD IN <= 41'b10111011000000000000000000000000000001001;
$vcdplusoff;

end

initial begin
    $monitor($time, ": IN=%b, OUT=%b, SYN=%b, ERR=%b, SGL=%b, DBL=%b", IN, OUT, SYN, ERR, SGL, DBL);
end

endmodule

