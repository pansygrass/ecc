`timescale 1 ns /100 ps

module dec_32_tb();

reg [38:0] IN;
wire [38:0] OUT;
wire [6:0] SYN;
wire ERR, SGL, DBL;

sec_ded_dec_top DUT0 (.IN(IN), .FINOUT(OUT), .SYN(SYN), .ERR(ERR), .SGL(SGL), .DBL(DBL));
initial begin

$vcdpluson;
    IN <= 32'd0;
    #`CLOCK_PERIOD IN <= 32'b000000000000000000000000000000000000000;
    #`CLOCK_PERIOD IN <= 32'b000011100000000000000000000000000000001;
    #`CLOCK_PERIOD IN <= 32'b000101100000000000000000000000000000010;
    #`CLOCK_PERIOD IN <= 32'b000110000000000000000000000000000000011;
    #`CLOCK_PERIOD IN <= 32'b001001100000000000000000000000000000100;
    #`CLOCK_PERIOD IN <= 32'b001010000000000000000000000000000000101;
    #`CLOCK_PERIOD IN <= 32'b001100000000000000000000000000000000110;
    #`CLOCK_PERIOD IN <= 32'b001111100000000000000000000000000000111;
    #`CLOCK_PERIOD IN <= 32'b010001100000000000000000000000000001000;
    #`CLOCK_PERIOD IN <= 32'b010010000000000000000000000000000001001;
$vcdplusoff;

end

initial begin
    $monitor($time, ": IN=%b, OUT=%b, ERR=%b, SGL=%b, DBL=%b", IN, OUT, ERR, SGL, DBL);
end

endmodule

