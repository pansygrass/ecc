VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO SRAM1R1W1024x32
  CLASS BLOCK ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 74.176 BY 63.232 ;
  SYMMETRY X Y R90 ;

  PIN CE1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 65.664 0.000 65.816 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 65.664 0.000 65.816 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 65.664 0.000 65.816 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 65.664 0.000 65.816 0.152 ;
    END
  END CE1

  PIN CSB1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 63.536 0.000 63.688 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 63.536 0.000 63.688 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 63.536 0.000 63.688 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 63.536 0.000 63.688 0.152 ;
    END
  END CSB1

  PIN OEB1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 61.408 0.000 61.560 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 61.408 0.000 61.560 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 61.408 0.000 61.560 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 61.408 0.000 61.560 0.152 ;
    END
  END OEB1

  PIN O1[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 59.280 0.000 59.432 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 59.280 0.000 59.432 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 59.280 0.000 59.432 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 59.280 0.000 59.432 0.152 ;
    END
  END O1[3]

  PIN O1[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 58.976 0.000 59.128 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 58.976 0.000 59.128 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 58.976 0.000 59.128 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 58.976 0.000 59.128 0.152 ;
    END
  END O1[2]

  PIN O1[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 58.672 0.000 58.824 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 58.672 0.000 58.824 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 58.672 0.000 58.824 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 58.672 0.000 58.824 0.152 ;
    END
  END O1[1]

  PIN O1[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 58.368 0.000 58.520 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 58.368 0.000 58.520 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 58.368 0.000 58.520 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 58.368 0.000 58.520 0.152 ;
    END
  END O1[0]

  PIN O1[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 56.240 0.000 56.392 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 56.240 0.000 56.392 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 56.240 0.000 56.392 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 56.240 0.000 56.392 0.152 ;
    END
  END O1[7]

  PIN O1[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 55.936 0.000 56.088 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 55.936 0.000 56.088 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 55.936 0.000 56.088 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 55.936 0.000 56.088 0.152 ;
    END
  END O1[6]

  PIN O1[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 55.632 0.000 55.784 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 55.632 0.000 55.784 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 55.632 0.000 55.784 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 55.632 0.000 55.784 0.152 ;
    END
  END O1[5]

  PIN O1[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 55.328 0.000 55.480 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 55.328 0.000 55.480 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 55.328 0.000 55.480 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 55.328 0.000 55.480 0.152 ;
    END
  END O1[4]

  PIN O1[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 53.200 0.000 53.352 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 53.200 0.000 53.352 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 53.200 0.000 53.352 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 53.200 0.000 53.352 0.152 ;
    END
  END O1[11]

  PIN O1[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 52.896 0.000 53.048 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 52.896 0.000 53.048 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 52.896 0.000 53.048 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 52.896 0.000 53.048 0.152 ;
    END
  END O1[10]

  PIN O1[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 52.592 0.000 52.744 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 52.592 0.000 52.744 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 52.592 0.000 52.744 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 52.592 0.000 52.744 0.152 ;
    END
  END O1[9]

  PIN O1[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 52.288 0.000 52.440 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 52.288 0.000 52.440 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 52.288 0.000 52.440 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 52.288 0.000 52.440 0.152 ;
    END
  END O1[8]

  PIN O1[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 50.160 0.000 50.312 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 50.160 0.000 50.312 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 50.160 0.000 50.312 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 50.160 0.000 50.312 0.152 ;
    END
  END O1[15]

  PIN O1[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 49.856 0.000 50.008 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 49.856 0.000 50.008 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 49.856 0.000 50.008 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 49.856 0.000 50.008 0.152 ;
    END
  END O1[14]

  PIN O1[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 49.552 0.000 49.704 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 49.552 0.000 49.704 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 49.552 0.000 49.704 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 49.552 0.000 49.704 0.152 ;
    END
  END O1[13]

  PIN O1[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 49.248 0.000 49.400 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 49.248 0.000 49.400 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 49.248 0.000 49.400 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 49.248 0.000 49.400 0.152 ;
    END
  END O1[12]

  PIN O1[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 47.120 0.000 47.272 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 47.120 0.000 47.272 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 47.120 0.000 47.272 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 47.120 0.000 47.272 0.152 ;
    END
  END O1[19]

  PIN O1[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 46.816 0.000 46.968 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 46.816 0.000 46.968 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 46.816 0.000 46.968 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 46.816 0.000 46.968 0.152 ;
    END
  END O1[18]

  PIN O1[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 46.512 0.000 46.664 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 46.512 0.000 46.664 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 46.512 0.000 46.664 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 46.512 0.000 46.664 0.152 ;
    END
  END O1[17]

  PIN O1[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 46.208 0.000 46.360 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 46.208 0.000 46.360 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 46.208 0.000 46.360 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 46.208 0.000 46.360 0.152 ;
    END
  END O1[16]

  PIN O1[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 44.080 0.000 44.232 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 44.080 0.000 44.232 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 44.080 0.000 44.232 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 44.080 0.000 44.232 0.152 ;
    END
  END O1[23]

  PIN O1[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 43.776 0.000 43.928 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 43.776 0.000 43.928 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 43.776 0.000 43.928 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 43.776 0.000 43.928 0.152 ;
    END
  END O1[22]

  PIN O1[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 43.472 0.000 43.624 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 43.472 0.000 43.624 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 43.472 0.000 43.624 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 43.472 0.000 43.624 0.152 ;
    END
  END O1[21]

  PIN O1[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 43.168 0.000 43.320 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 43.168 0.000 43.320 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 43.168 0.000 43.320 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 43.168 0.000 43.320 0.152 ;
    END
  END O1[20]

  PIN O1[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 41.040 0.000 41.192 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 41.040 0.000 41.192 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 41.040 0.000 41.192 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 41.040 0.000 41.192 0.152 ;
    END
  END O1[27]

  PIN O1[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 40.736 0.000 40.888 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 40.736 0.000 40.888 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 40.736 0.000 40.888 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 40.736 0.000 40.888 0.152 ;
    END
  END O1[26]

  PIN O1[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 40.432 0.000 40.584 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 40.432 0.000 40.584 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 40.432 0.000 40.584 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 40.432 0.000 40.584 0.152 ;
    END
  END O1[25]

  PIN O1[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 40.128 0.000 40.280 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 40.128 0.000 40.280 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 40.128 0.000 40.280 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 40.128 0.000 40.280 0.152 ;
    END
  END O1[24]

  PIN O1[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 38.000 0.000 38.152 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 38.000 0.000 38.152 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 38.000 0.000 38.152 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 38.000 0.000 38.152 0.152 ;
    END
  END O1[31]

  PIN O1[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 37.696 0.000 37.848 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 37.696 0.000 37.848 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 37.696 0.000 37.848 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 37.696 0.000 37.848 0.152 ;
    END
  END O1[30]

  PIN O1[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 37.392 0.000 37.544 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 37.392 0.000 37.544 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 37.392 0.000 37.544 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 37.392 0.000 37.544 0.152 ;
    END
  END O1[29]

  PIN O1[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 37.088 0.000 37.240 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 37.088 0.000 37.240 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 37.088 0.000 37.240 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 37.088 0.000 37.240 0.152 ;
    END
  END O1[28]

  PIN A1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 74.024 55.328 74.176 55.480 ;
    END
    PORT
      LAYER M3 ;
        RECT 74.024 55.328 74.176 55.480 ;
    END
    PORT
      LAYER M4 ;
        RECT 74.024 55.328 74.176 55.480 ;
    END
    PORT
      LAYER M5 ;
        RECT 74.024 55.328 74.176 55.480 ;
    END
  END A1[0]

  PIN A1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 74.024 51.680 74.176 51.832 ;
    END
    PORT
      LAYER M3 ;
        RECT 74.024 51.680 74.176 51.832 ;
    END
    PORT
      LAYER M4 ;
        RECT 74.024 51.680 74.176 51.832 ;
    END
    PORT
      LAYER M5 ;
        RECT 74.024 51.680 74.176 51.832 ;
    END
  END A1[1]

  PIN A1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 74.024 48.032 74.176 48.184 ;
    END
    PORT
      LAYER M3 ;
        RECT 74.024 48.032 74.176 48.184 ;
    END
    PORT
      LAYER M4 ;
        RECT 74.024 48.032 74.176 48.184 ;
    END
    PORT
      LAYER M5 ;
        RECT 74.024 48.032 74.176 48.184 ;
    END
  END A1[2]

  PIN A1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 74.024 44.384 74.176 44.536 ;
    END
    PORT
      LAYER M3 ;
        RECT 74.024 44.384 74.176 44.536 ;
    END
    PORT
      LAYER M4 ;
        RECT 74.024 44.384 74.176 44.536 ;
    END
    PORT
      LAYER M5 ;
        RECT 74.024 44.384 74.176 44.536 ;
    END
  END A1[3]

  PIN A1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 74.024 40.736 74.176 40.888 ;
    END
    PORT
      LAYER M3 ;
        RECT 74.024 40.736 74.176 40.888 ;
    END
    PORT
      LAYER M4 ;
        RECT 74.024 40.736 74.176 40.888 ;
    END
    PORT
      LAYER M5 ;
        RECT 74.024 40.736 74.176 40.888 ;
    END
  END A1[4]

  PIN A1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 74.024 37.088 74.176 37.240 ;
    END
    PORT
      LAYER M3 ;
        RECT 74.024 37.088 74.176 37.240 ;
    END
    PORT
      LAYER M4 ;
        RECT 74.024 37.088 74.176 37.240 ;
    END
    PORT
      LAYER M5 ;
        RECT 74.024 37.088 74.176 37.240 ;
    END
  END A1[5]

  PIN A1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 74.024 33.440 74.176 33.592 ;
    END
    PORT
      LAYER M3 ;
        RECT 74.024 33.440 74.176 33.592 ;
    END
    PORT
      LAYER M4 ;
        RECT 74.024 33.440 74.176 33.592 ;
    END
    PORT
      LAYER M5 ;
        RECT 74.024 33.440 74.176 33.592 ;
    END
  END A1[6]

  PIN A1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 74.024 29.792 74.176 29.944 ;
    END
    PORT
      LAYER M3 ;
        RECT 74.024 29.792 74.176 29.944 ;
    END
    PORT
      LAYER M4 ;
        RECT 74.024 29.792 74.176 29.944 ;
    END
    PORT
      LAYER M5 ;
        RECT 74.024 29.792 74.176 29.944 ;
    END
  END A1[7]

  PIN CE2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8.512 0.000 8.664 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 8.512 0.000 8.664 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 8.512 0.000 8.664 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 8.512 0.000 8.664 0.152 ;
    END
  END CE2

  PIN CSB2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10.640 0.000 10.792 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 10.640 0.000 10.792 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 10.640 0.000 10.792 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 10.640 0.000 10.792 0.152 ;
    END
  END CSB2

  PIN I2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12.768 0.000 12.920 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 12.768 0.000 12.920 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 12.768 0.000 12.920 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 12.768 0.000 12.920 0.152 ;
    END
  END I2[0]

  PIN I2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13.072 0.000 13.224 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 13.072 0.000 13.224 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 13.072 0.000 13.224 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 13.072 0.000 13.224 0.152 ;
    END
  END I2[1]

  PIN I2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13.376 0.000 13.528 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 13.376 0.000 13.528 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 13.376 0.000 13.528 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 13.376 0.000 13.528 0.152 ;
    END
  END I2[2]

  PIN I2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13.680 0.000 13.832 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 13.680 0.000 13.832 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 13.680 0.000 13.832 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 13.680 0.000 13.832 0.152 ;
    END
  END I2[3]

  PIN I2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15.808 0.000 15.960 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 15.808 0.000 15.960 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 15.808 0.000 15.960 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 15.808 0.000 15.960 0.152 ;
    END
  END I2[4]

  PIN I2[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16.112 0.000 16.264 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 16.112 0.000 16.264 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 16.112 0.000 16.264 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 16.112 0.000 16.264 0.152 ;
    END
  END I2[5]

  PIN I2[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16.416 0.000 16.568 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 16.416 0.000 16.568 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 16.416 0.000 16.568 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 16.416 0.000 16.568 0.152 ;
    END
  END I2[6]

  PIN I2[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16.720 0.000 16.872 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 16.720 0.000 16.872 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 16.720 0.000 16.872 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 16.720 0.000 16.872 0.152 ;
    END
  END I2[7]

  PIN I2[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18.848 0.000 19.000 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 18.848 0.000 19.000 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 18.848 0.000 19.000 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 18.848 0.000 19.000 0.152 ;
    END
  END I2[8]

  PIN I2[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 19.152 0.000 19.304 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 19.152 0.000 19.304 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 19.152 0.000 19.304 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 19.152 0.000 19.304 0.152 ;
    END
  END I2[9]

  PIN I2[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 19.456 0.000 19.608 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 19.456 0.000 19.608 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 19.456 0.000 19.608 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 19.456 0.000 19.608 0.152 ;
    END
  END I2[10]

  PIN I2[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 19.760 0.000 19.912 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 19.760 0.000 19.912 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 19.760 0.000 19.912 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 19.760 0.000 19.912 0.152 ;
    END
  END I2[11]

  PIN I2[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 21.888 0.000 22.040 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 21.888 0.000 22.040 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 21.888 0.000 22.040 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 21.888 0.000 22.040 0.152 ;
    END
  END I2[12]

  PIN I2[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 22.192 0.000 22.344 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 22.192 0.000 22.344 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 22.192 0.000 22.344 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 22.192 0.000 22.344 0.152 ;
    END
  END I2[13]

  PIN I2[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 22.496 0.000 22.648 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 22.496 0.000 22.648 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 22.496 0.000 22.648 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 22.496 0.000 22.648 0.152 ;
    END
  END I2[14]

  PIN I2[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 22.800 0.000 22.952 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 22.800 0.000 22.952 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 22.800 0.000 22.952 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 22.800 0.000 22.952 0.152 ;
    END
  END I2[15]

  PIN I2[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 24.928 0.000 25.080 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 24.928 0.000 25.080 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 24.928 0.000 25.080 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 24.928 0.000 25.080 0.152 ;
    END
  END I2[16]

  PIN I2[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 25.232 0.000 25.384 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 25.232 0.000 25.384 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 25.232 0.000 25.384 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 25.232 0.000 25.384 0.152 ;
    END
  END I2[17]

  PIN I2[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 25.536 0.000 25.688 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 25.536 0.000 25.688 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 25.536 0.000 25.688 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 25.536 0.000 25.688 0.152 ;
    END
  END I2[18]

  PIN I2[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 25.840 0.000 25.992 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 25.840 0.000 25.992 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 25.840 0.000 25.992 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 25.840 0.000 25.992 0.152 ;
    END
  END I2[19]

  PIN I2[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 27.968 0.000 28.120 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 27.968 0.000 28.120 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 27.968 0.000 28.120 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 27.968 0.000 28.120 0.152 ;
    END
  END I2[20]

  PIN I2[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 28.272 0.000 28.424 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 28.272 0.000 28.424 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 28.272 0.000 28.424 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 28.272 0.000 28.424 0.152 ;
    END
  END I2[21]

  PIN I2[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 28.576 0.000 28.728 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 28.576 0.000 28.728 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 28.576 0.000 28.728 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 28.576 0.000 28.728 0.152 ;
    END
  END I2[22]

  PIN I2[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 28.880 0.000 29.032 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 28.880 0.000 29.032 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 28.880 0.000 29.032 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 28.880 0.000 29.032 0.152 ;
    END
  END I2[23]

  PIN I2[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 31.008 0.000 31.160 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 31.008 0.000 31.160 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 31.008 0.000 31.160 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 31.008 0.000 31.160 0.152 ;
    END
  END I2[24]

  PIN I2[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 31.312 0.000 31.464 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 31.312 0.000 31.464 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 31.312 0.000 31.464 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 31.312 0.000 31.464 0.152 ;
    END
  END I2[25]

  PIN I2[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 31.616 0.000 31.768 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 31.616 0.000 31.768 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 31.616 0.000 31.768 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 31.616 0.000 31.768 0.152 ;
    END
  END I2[26]

  PIN I2[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 31.920 0.000 32.072 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 31.920 0.000 32.072 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 31.920 0.000 32.072 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 31.920 0.000 32.072 0.152 ;
    END
  END I2[27]

  PIN I2[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 34.048 0.000 34.200 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 34.048 0.000 34.200 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 34.048 0.000 34.200 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 34.048 0.000 34.200 0.152 ;
    END
  END I2[28]

  PIN I2[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 34.352 0.000 34.504 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 34.352 0.000 34.504 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 34.352 0.000 34.504 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 34.352 0.000 34.504 0.152 ;
    END
  END I2[29]

  PIN I2[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 34.656 0.000 34.808 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 34.656 0.000 34.808 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 34.656 0.000 34.808 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 34.656 0.000 34.808 0.152 ;
    END
  END I2[30]

  PIN I2[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 34.960 0.000 35.112 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 34.960 0.000 35.112 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 34.960 0.000 35.112 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 34.960 0.000 35.112 0.152 ;
    END
  END I2[31]

  PIN A2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.000 55.328 0.152 55.480 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.000 55.328 0.152 55.480 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.000 55.328 0.152 55.480 ;
    END
    PORT
      LAYER M5 ;
        RECT 0.000 55.328 0.152 55.480 ;
    END
  END A2[0]

  PIN A2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.000 51.680 0.152 51.832 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.000 51.680 0.152 51.832 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.000 51.680 0.152 51.832 ;
    END
    PORT
      LAYER M5 ;
        RECT 0.000 51.680 0.152 51.832 ;
    END
  END A2[1]

  PIN A2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.000 48.032 0.152 48.184 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.000 48.032 0.152 48.184 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.000 48.032 0.152 48.184 ;
    END
    PORT
      LAYER M5 ;
        RECT 0.000 48.032 0.152 48.184 ;
    END
  END A2[2]

  PIN A2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.000 44.384 0.152 44.536 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.000 44.384 0.152 44.536 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.000 44.384 0.152 44.536 ;
    END
    PORT
      LAYER M5 ;
        RECT 0.000 44.384 0.152 44.536 ;
    END
  END A2[3]

  PIN A2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.000 40.736 0.152 40.888 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.000 40.736 0.152 40.888 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.000 40.736 0.152 40.888 ;
    END
    PORT
      LAYER M5 ;
        RECT 0.000 40.736 0.152 40.888 ;
    END
  END A2[4]

  PIN A2[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.000 37.088 0.152 37.240 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.000 37.088 0.152 37.240 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.000 37.088 0.152 37.240 ;
    END
    PORT
      LAYER M5 ;
        RECT 0.000 37.088 0.152 37.240 ;
    END
  END A2[5]

  PIN A2[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.000 33.440 0.152 33.592 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.000 33.440 0.152 33.592 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.000 33.440 0.152 33.592 ;
    END
    PORT
      LAYER M5 ;
        RECT 0.000 33.440 0.152 33.592 ;
    END
  END A2[6]

  PIN A2[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.000 29.792 0.152 29.944 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.000 29.792 0.152 29.944 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.000 29.792 0.152 29.944 ;
    END
    PORT
      LAYER M5 ;
        RECT 0.000 29.792 0.152 29.944 ;
    END
  END A2[7]

  PIN WEB2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.000 15.808 0.152 15.960 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.000 15.808 0.152 15.960 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.000 15.808 0.152 15.960 ;
    END
    PORT
      LAYER M5 ;
        RECT 0.000 15.808 0.152 15.960 ;
    END
  END WEB2

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M2 ;
        RECT 5.195 61.232 7.195 63.232 ;
    END
    PORT
      LAYER M3 ;
        RECT 5.195 61.232 7.195 63.232 ;
    END
    PORT
      LAYER M5 ;
        RECT 5.195 61.232 7.195 63.232 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M2 ;
        RECT 7.915 61.232 9.915 63.232 ;
    END
    PORT
      LAYER M3 ;
        RECT 7.915 61.232 9.915 63.232 ;
    END
    PORT
      LAYER M5 ;
        RECT 7.915 61.232 9.915 63.232 ;
    END
  END VSS

  OBS
    LAYER M2 ;
      RECT 65.968 0.000 74.176 0.304 ;
      RECT 63.840 0.000 65.512 0.304 ;
      RECT 61.712 0.000 63.384 0.304 ;
      RECT 59.584 0.000 61.256 0.304 ;
      RECT 56.544 0.000 58.216 0.304 ;
      RECT 53.504 0.000 55.176 0.304 ;
      RECT 50.464 0.000 52.136 0.304 ;
      RECT 47.424 0.000 49.096 0.304 ;
      RECT 44.384 0.000 46.056 0.304 ;
      RECT 41.344 0.000 43.016 0.304 ;
      RECT 38.304 0.000 39.976 0.304 ;
      RECT 73.872 55.632 74.176 61.080 ;
      RECT 73.872 51.984 74.176 55.176 ;
      RECT 73.872 48.336 74.176 51.528 ;
      RECT 73.872 44.688 74.176 47.880 ;
      RECT 73.872 41.040 74.176 44.232 ;
      RECT 73.872 37.392 74.176 40.584 ;
      RECT 73.872 33.744 74.176 36.936 ;
      RECT 73.872 30.096 74.176 33.288 ;
      RECT 73.872 16.112 74.176 29.640 ;
      RECT 73.872 0.304 74.176 15.656 ;
      RECT 0.000 0.000 8.360 0.304 ;
      RECT 8.816 0.000 10.488 0.304 ;
      RECT 10.944 0.000 12.616 0.304 ;
      RECT 13.984 0.000 15.656 0.304 ;
      RECT 17.024 0.000 18.696 0.304 ;
      RECT 20.064 0.000 21.736 0.304 ;
      RECT 23.104 0.000 24.776 0.304 ;
      RECT 26.144 0.000 27.816 0.304 ;
      RECT 29.184 0.000 30.856 0.304 ;
      RECT 32.224 0.000 33.896 0.304 ;
      RECT 35.264 0.000 36.936 0.304 ;
      RECT 0.000 55.632 0.304 61.080 ;
      RECT 0.000 51.984 0.304 55.176 ;
      RECT 0.000 48.336 0.304 51.528 ;
      RECT 0.000 44.688 0.304 47.880 ;
      RECT 0.000 41.040 0.304 44.232 ;
      RECT 0.000 37.392 0.304 40.584 ;
      RECT 0.000 33.744 0.304 36.936 ;
      RECT 0.000 30.096 0.304 33.288 ;
      RECT 0.000 16.112 0.304 29.640 ;
      RECT 0.000 0.304 0.304 15.656 ;
      RECT 0.000 61.080 5.043 63.232 ;
      RECT 7.355 61.080 7.763 63.232 ;
      RECT 10.067 61.080 74.176 63.232 ;
      RECT 0.304 0.304 73.872 61.080 ;
    LAYER M3 ;
      RECT 65.968 0.000 74.176 0.304 ;
      RECT 63.840 0.000 65.512 0.304 ;
      RECT 61.712 0.000 63.384 0.304 ;
      RECT 59.584 0.000 61.256 0.304 ;
      RECT 56.544 0.000 58.216 0.304 ;
      RECT 53.504 0.000 55.176 0.304 ;
      RECT 50.464 0.000 52.136 0.304 ;
      RECT 47.424 0.000 49.096 0.304 ;
      RECT 44.384 0.000 46.056 0.304 ;
      RECT 41.344 0.000 43.016 0.304 ;
      RECT 38.304 0.000 39.976 0.304 ;
      RECT 73.872 55.632 74.176 61.080 ;
      RECT 73.872 51.984 74.176 55.176 ;
      RECT 73.872 48.336 74.176 51.528 ;
      RECT 73.872 44.688 74.176 47.880 ;
      RECT 73.872 41.040 74.176 44.232 ;
      RECT 73.872 37.392 74.176 40.584 ;
      RECT 73.872 33.744 74.176 36.936 ;
      RECT 73.872 30.096 74.176 33.288 ;
      RECT 73.872 16.112 74.176 29.640 ;
      RECT 73.872 0.304 74.176 15.656 ;
      RECT 0.000 0.000 8.360 0.304 ;
      RECT 8.816 0.000 10.488 0.304 ;
      RECT 10.944 0.000 12.616 0.304 ;
      RECT 13.984 0.000 15.656 0.304 ;
      RECT 17.024 0.000 18.696 0.304 ;
      RECT 20.064 0.000 21.736 0.304 ;
      RECT 23.104 0.000 24.776 0.304 ;
      RECT 26.144 0.000 27.816 0.304 ;
      RECT 29.184 0.000 30.856 0.304 ;
      RECT 32.224 0.000 33.896 0.304 ;
      RECT 35.264 0.000 36.936 0.304 ;
      RECT 0.000 55.632 0.304 61.080 ;
      RECT 0.000 51.984 0.304 55.176 ;
      RECT 0.000 48.336 0.304 51.528 ;
      RECT 0.000 44.688 0.304 47.880 ;
      RECT 0.000 41.040 0.304 44.232 ;
      RECT 0.000 37.392 0.304 40.584 ;
      RECT 0.000 33.744 0.304 36.936 ;
      RECT 0.000 30.096 0.304 33.288 ;
      RECT 0.000 16.112 0.304 29.640 ;
      RECT 0.000 0.304 0.304 15.656 ;
      RECT 0.000 61.080 5.043 63.232 ;
      RECT 7.355 61.080 7.763 63.232 ;
      RECT 10.067 61.080 74.176 63.232 ;
      RECT 0.304 0.304 73.872 61.080 ;
    LAYER M4 ;
      RECT 65.968 0.000 74.176 0.304 ;
      RECT 63.840 0.000 65.512 0.304 ;
      RECT 61.712 0.000 63.384 0.304 ;
      RECT 59.584 0.000 61.256 0.304 ;
      RECT 56.544 0.000 58.216 0.304 ;
      RECT 53.504 0.000 55.176 0.304 ;
      RECT 50.464 0.000 52.136 0.304 ;
      RECT 47.424 0.000 49.096 0.304 ;
      RECT 44.384 0.000 46.056 0.304 ;
      RECT 41.344 0.000 43.016 0.304 ;
      RECT 38.304 0.000 39.976 0.304 ;
      RECT 73.872 55.632 74.176 61.080 ;
      RECT 73.872 51.984 74.176 55.176 ;
      RECT 73.872 48.336 74.176 51.528 ;
      RECT 73.872 44.688 74.176 47.880 ;
      RECT 73.872 41.040 74.176 44.232 ;
      RECT 73.872 37.392 74.176 40.584 ;
      RECT 73.872 33.744 74.176 36.936 ;
      RECT 73.872 30.096 74.176 33.288 ;
      RECT 73.872 16.112 74.176 29.640 ;
      RECT 73.872 0.304 74.176 15.656 ;
      RECT 0.000 0.000 8.360 0.304 ;
      RECT 8.816 0.000 10.488 0.304 ;
      RECT 10.944 0.000 12.616 0.304 ;
      RECT 13.984 0.000 15.656 0.304 ;
      RECT 17.024 0.000 18.696 0.304 ;
      RECT 20.064 0.000 21.736 0.304 ;
      RECT 23.104 0.000 24.776 0.304 ;
      RECT 26.144 0.000 27.816 0.304 ;
      RECT 29.184 0.000 30.856 0.304 ;
      RECT 32.224 0.000 33.896 0.304 ;
      RECT 35.264 0.000 36.936 0.304 ;
      RECT 0.000 55.632 0.304 61.080 ;
      RECT 0.000 51.984 0.304 55.176 ;
      RECT 0.000 48.336 0.304 51.528 ;
      RECT 0.000 44.688 0.304 47.880 ;
      RECT 0.000 41.040 0.304 44.232 ;
      RECT 0.000 37.392 0.304 40.584 ;
      RECT 0.000 33.744 0.304 36.936 ;
      RECT 0.000 30.096 0.304 33.288 ;
      RECT 0.000 16.112 0.304 29.640 ;
      RECT 0.000 0.304 0.304 15.656 ;
      RECT 0.000 61.080 5.043 63.232 ;
      RECT 7.355 61.080 7.763 63.232 ;
      RECT 10.067 61.080 74.176 63.232 ;
      RECT 0.304 0.304 73.872 61.080 ;
    LAYER M5 ;
      RECT 65.968 0.000 74.176 0.304 ;
      RECT 63.840 0.000 65.512 0.304 ;
      RECT 61.712 0.000 63.384 0.304 ;
      RECT 59.584 0.000 61.256 0.304 ;
      RECT 56.544 0.000 58.216 0.304 ;
      RECT 53.504 0.000 55.176 0.304 ;
      RECT 50.464 0.000 52.136 0.304 ;
      RECT 47.424 0.000 49.096 0.304 ;
      RECT 44.384 0.000 46.056 0.304 ;
      RECT 41.344 0.000 43.016 0.304 ;
      RECT 38.304 0.000 39.976 0.304 ;
      RECT 73.872 55.632 74.176 61.080 ;
      RECT 73.872 51.984 74.176 55.176 ;
      RECT 73.872 48.336 74.176 51.528 ;
      RECT 73.872 44.688 74.176 47.880 ;
      RECT 73.872 41.040 74.176 44.232 ;
      RECT 73.872 37.392 74.176 40.584 ;
      RECT 73.872 33.744 74.176 36.936 ;
      RECT 73.872 30.096 74.176 33.288 ;
      RECT 73.872 16.112 74.176 29.640 ;
      RECT 73.872 0.304 74.176 15.656 ;
      RECT 0.000 0.000 8.360 0.304 ;
      RECT 8.816 0.000 10.488 0.304 ;
      RECT 10.944 0.000 12.616 0.304 ;
      RECT 13.984 0.000 15.656 0.304 ;
      RECT 17.024 0.000 18.696 0.304 ;
      RECT 20.064 0.000 21.736 0.304 ;
      RECT 23.104 0.000 24.776 0.304 ;
      RECT 26.144 0.000 27.816 0.304 ;
      RECT 29.184 0.000 30.856 0.304 ;
      RECT 32.224 0.000 33.896 0.304 ;
      RECT 35.264 0.000 36.936 0.304 ;
      RECT 0.000 55.632 0.304 61.080 ;
      RECT 0.000 51.984 0.304 55.176 ;
      RECT 0.000 48.336 0.304 51.528 ;
      RECT 0.000 44.688 0.304 47.880 ;
      RECT 0.000 41.040 0.304 44.232 ;
      RECT 0.000 37.392 0.304 40.584 ;
      RECT 0.000 33.744 0.304 36.936 ;
      RECT 0.000 30.096 0.304 33.288 ;
      RECT 0.000 16.112 0.304 29.640 ;
      RECT 0.000 0.304 0.304 15.656 ;
      RECT 0.000 61.080 5.043 63.232 ;
      RECT 7.355 61.080 7.763 63.232 ;
      RECT 10.067 61.080 74.176 63.232 ;
      RECT 0.304 0.304 73.872 61.080 ;
  END

END SRAM1R1W1024x32

END LIBRARY
