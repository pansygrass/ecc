//
// decoder for Hsiao 128 bit SEC-DED
//
// Authors: Joseph Crowe and Matt Markwell
//


module corrector (input [126:0] IN, 
    input [13:0] SYN,
    output reg [126:0] OUT
);

reg [126:0] LOC;

    always @(*) begin
        case(SYN)

14'h0377 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001; // S (0x00000000000000000000000000000001) 
14'h0599 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011; // D (0x00000000000000000000000000000003) 
14'h0eab : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101; // D (0x00000000000000000000000000000005) 
14'h18cf : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001; // D (0x00000000000000000000000000000009) 
14'h3407 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001; // D (0x00000000000000000000000000000011) 
14'h2ee0 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100001; // D (0x00000000000000000000000000000021) 
14'h1b2e : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000001; // D (0x00000000000000000000000000000041) 
14'h33c5 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000001; // D (0x00000000000000000000000000000081) 
14'h2164 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000001; // D (0x00000000000000000000000000000101) 
14'h0426 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000001; // D (0x00000000000000000000000000000201) 
14'h0dd5 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000001; // D (0x00000000000000000000000000000401) 
14'h1e33 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000001; // D (0x00000000000000000000000000000801) 
14'h39ff : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000001; // D (0x00000000000000000000000000001001) 
14'h3510 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000001; // D (0x00000000000000000000000000002001) 
14'h2cce : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000001; // D (0x00000000000000000000000000004001) 
14'h1f72 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000001; // D (0x00000000000000000000000000008001) 
14'h3b7d : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001; // D (0x00000000000000000000000000010001) 
14'h3014 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000001; // D (0x00000000000000000000000000020001) 
14'h26c6 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000001; // D (0x00000000000000000000000000040001) 
14'h0b62 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000001; // D (0x00000000000000000000000000080001) 
14'h135d : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000001; // D (0x00000000000000000000000000100001) 
14'h2323 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000001; // D (0x00000000000000000000000000200001) 
14'h00a8 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000001; // D (0x00000000000000000000000000400001) 
14'h04c9 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000001; // D (0x00000000000000000000000000800001) 
14'h0c0b : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000001; // D (0x00000000000000000000000001000001) 
14'h1d8f : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000001; // D (0x00000000000000000000000002000001) 
14'h3e87 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000001; // D (0x00000000000000000000000004000001) 
14'h3be0 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000001; // D (0x00000000000000000000000008000001) 
14'h312e : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000001; // D (0x00000000000000000000000010000001) 
14'h24b2 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000001; // D (0x00000000000000000000000020000001) 
14'h0f8a : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000001; // D (0x00000000000000000000000040000001) 
14'h1a8d : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000001; // D (0x00000000000000000000000080000001) 
14'h3083 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000001; // D (0x00000000000000000000000100000001) 
14'h27e8 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000001; // D (0x00000000000000000000000200000001) 
14'h093e : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000001; // D (0x00000000000000000000000400000001) 
14'h17e5 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000001; // D (0x00000000000000000000000800000001) 
14'h2a53 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000001; // D (0x00000000000000000000001000000001) 
14'h1248 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000001; // D (0x00000000000000000000002000000001) 
14'h2109 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000001; // D (0x00000000000000000000004000000001) 
14'h04fc : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000001; // D (0x00000000000000000000008000000001) 
14'h0c61 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000001; // D (0x00000000000000000000010000000001) 
14'h1d5b : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000001; // D (0x00000000000000000000020000000001) 
14'h3f2f : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000001; // D (0x00000000000000000000040000000001) 
14'h38b0 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000001; // D (0x00000000000000000000080000000001) 
14'h378e : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000001; // D (0x00000000000000000000100000000001) 
14'h29f2 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000001; // D (0x00000000000000000000200000000001) 
14'h150a : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000001; // D (0x00000000000000000000400000000001) 
14'h2f8d : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000001; // D (0x00000000000000000000800000000001) 
14'h19f4 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000001; // D (0x00000000000000000001000000000001) 
14'h3671 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000001; // D (0x00000000000000000002000000000001) 
14'h2a0c : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000001; // D (0x00000000000000000004000000000001) 
14'h12f6 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000001; // D (0x00000000000000000008000000000001) 
14'h2075 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000001; // D (0x00000000000000000010000000000001) 
14'h0604 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000001; // D (0x00000000000000000020000000000001) 
14'h0991 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000001; // D (0x00000000000000000040000000000001) 
14'h16bb : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000001; // D (0x00000000000000000080000000000001) 
14'h28ef : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000001; // D (0x00000000000000000100000000000001) 
14'h1730 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000001; // D (0x00000000000000000200000000000001) 
14'h2bf9 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000001; // D (0x00000000000000000400000000000001) 
14'h111c : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000001; // D (0x00000000000000000800000000000001) 
14'h27a1 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000001; // D (0x00000000000000001000000000000001) 
14'h09ac : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000001; // D (0x00000000000000002000000000000001) 
14'h16c1 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000001; // D (0x00000000000000004000000000000001) 
14'h281b : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000001; // D (0x00000000000000008000000000000001) 
14'h16d8 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000001; // D (0x00000000000000010000000000000001) 
14'h2829 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000001; // D (0x00000000000000020000000000000001) 
14'h16bc : LOC =         127'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000001; // D (0x00000000000000040000000000000001) 
14'h28e1 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000001; // D (0x00000000000000080000000000000001) 
14'h172c : LOC =         127'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000001; // D (0x00000000000000100000000000000001) 
14'h2bc1 : LOC =         127'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000001; // D (0x00000000000000200000000000000001) 
14'h116c : LOC =         127'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000001; // D (0x00000000000000400000000000000001) 
14'h2741 : LOC =         127'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000001; // D (0x00000000000000800000000000000001) 
14'h086c : LOC =         127'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000001; // D (0x00000000000001000000000000000001) 
14'h1541 : LOC =         127'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000001; // D (0x00000000000002000000000000000001) 
14'h2f1b : LOC =         127'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000001; // D (0x00000000000004000000000000000001) 
14'h18d8 : LOC =         127'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000001; // D (0x00000000000008000000000000000001) 
14'h3429 : LOC =         127'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000001; // D (0x00000000000010000000000000000001) 
14'h2ebc : LOC =         127'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000001; // D (0x00000000000020000000000000000001) 
14'h1b96 : LOC =         127'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000001; // D (0x00000000000040000000000000000001) 
14'h32b5 : LOC =         127'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000001; // D (0x00000000000080000000000000000001) 
14'h2384 : LOC =         127'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000001; // D (0x00000000000100000000000000000001) 
14'h01e6 : LOC =         127'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000001; // D (0x00000000000200000000000000000001) 
14'h0655 : LOC =         127'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000001; // D (0x00000000000400000000000000000001) 
14'h0933 : LOC =         127'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000001; // D (0x00000000000800000000000000000001) 
14'h17ff : LOC =         127'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000001; // D (0x00000000001000000000000000000001) 
14'h2a67 : LOC =         127'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000001; // D (0x00000000002000000000000000000001) 
14'h1220 : LOC =         127'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000001; // D (0x00000000004000000000000000000001) 
14'h21d9 : LOC =         127'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000001; // D (0x00000000008000000000000000000001) 
14'h055c : LOC =         127'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000001; // D (0x00000000010000000000000000000001) 
14'h0f21 : LOC =         127'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000001; // D (0x00000000020000000000000000000001) 
14'h1bdb : LOC =         127'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001; // D (0x00000000040000000000000000000001) 
14'h322f : LOC =         127'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001; // D (0x00000000080000000000000000000001) 
14'h22b0 : LOC =         127'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001; // D (0x00000000100000000000000000000001) 
14'h038e : LOC =         127'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001; // D (0x00000000200000000000000000000001) 
14'h0285 : LOC =         127'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001; // D (0x00000000400000000000000000000001) 
14'h0093 : LOC =         127'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001; // D (0x00000000800000000000000000000001) 
14'h04bf : LOC =         127'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001; // D (0x00000001000000000000000000000001) 
14'h0ce7 : LOC =         127'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001; // D (0x00000002000000000000000000000001) 
14'h1c57 : LOC =         127'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001; // D (0x00000004000000000000000000000001) 
14'h3d37 : LOC =         127'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001; // D (0x00000008000000000000000000000001) 
14'h3c80 : LOC =         127'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001; // D (0x00000010000000000000000000000001) 
14'h3fee : LOC =         127'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001; // D (0x00000020000000000000000000000001) 
14'h3932 : LOC =         127'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001; // D (0x00000040000000000000000000000001) 
14'h348a : LOC =         127'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001; // D (0x00000080000000000000000000000001) 
14'h2ffa : LOC =         127'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001; // D (0x00000100000000000000000000000001) 
14'h191a : LOC =         127'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001; // D (0x00000200000000000000000000000001) 
14'h37ad : LOC =         127'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001; // D (0x00000400000000000000000000000001) 
14'h29b4 : LOC =         127'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001; // D (0x00000800000000000000000000000001) 
14'h1586 : LOC =         127'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001; // D (0x00001000000000000000000000000001) 
14'h2e95 : LOC =         127'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001; // D (0x00002000000000000000000000000001) 
14'h1bc4 : LOC =         127'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001; // D (0x00004000000000000000000000000001) 
14'h3211 : LOC =         127'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001; // D (0x00008000000000000000000000000001) 
14'h22cc : LOC =         127'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001; // D (0x00010000000000000000000000000001) 
14'h0376 : LOC =         127'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001; // D (0x00020000000000000000000000000001) 
14'h0375 : LOC =         127'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001; // D (0x00040000000000000000000000000001) 
14'h0373 : LOC =         127'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001; // D (0x00080000000000000000000000000001) 
14'h037f : LOC =         127'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001; // D (0x00100000000000000000000000000001) 
14'h0367 : LOC =         127'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001; // D (0x00200000000000000000000000000001) 
14'h0357 : LOC =         127'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001; // D (0x00400000000000000000000000000001) 
14'h0337 : LOC =         127'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001; // D (0x00800000000000000000000000000001) 
14'h03f7 : LOC =         127'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001; // D (0x01000000000000000000000000000001) 
14'h0277 : LOC =         127'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001; // D (0x02000000000000000000000000000001) 
14'h0177 : LOC =         127'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001; // D (0x04000000000000000000000000000001) 
14'h0777 : LOC =         127'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001; // D (0x08000000000000000000000000000001) 
14'h0b77 : LOC =         127'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001; // D (0x10000000000000000000000000000001) 
14'h1377 : LOC =         127'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001; // D (0x20000000000000000000000000000001) 
14'h2377 : LOC =         127'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001; // D (0x40000000000000000000000000000001) 
14'h06ee : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010; // S (0x00000000000000000000000000000002) 
14'h0b32 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110; // D (0x00000000000000000000000000000006) 
14'h1d56 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010; // D (0x0000000000000000000000000000000a) 
14'h319e : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010; // D (0x00000000000000000000000000000012) 
14'h2b79 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010; // D (0x00000000000000000000000000000022) 
14'h1eb7 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000010; // D (0x00000000000000000000000000000042) 
14'h365c : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000010; // D (0x00000000000000000000000000000082) 
14'h24fd : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000010; // D (0x00000000000000000000000000000102) 
14'h01bf : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000010; // D (0x00000000000000000000000000000202) 
14'h084c : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000010; // D (0x00000000000000000000000000000402) 
14'h1baa : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000010; // D (0x00000000000000000000000000000802) 
14'h3c66 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000010; // D (0x00000000000000000000000000001002) 
14'h3089 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000010; // D (0x00000000000000000000000000002002) 
14'h2957 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000010; // D (0x00000000000000000000000000004002) 
14'h1aeb : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000010; // D (0x00000000000000000000000000008002) 
14'h3ee4 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000010; // D (0x00000000000000000000000000010002) 
14'h358d : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000010; // D (0x00000000000000000000000000020002) 
14'h235f : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000010; // D (0x00000000000000000000000000040002) 
14'h0efb : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000010; // D (0x00000000000000000000000000080002) 
14'h16c4 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000010; // D (0x00000000000000000000000000100002) 
14'h26ba : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000010; // D (0x00000000000000000000000000200002) 
14'h0531 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000010; // D (0x00000000000000000000000000400002) 
14'h0150 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000010; // D (0x00000000000000000000000000800002) 
14'h0992 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000010; // D (0x00000000000000000000000001000002) 
14'h1816 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000010; // D (0x00000000000000000000000002000002) 
14'h3b1e : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000010; // D (0x00000000000000000000000004000002) 
14'h3e79 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000010; // D (0x00000000000000000000000008000002) 
14'h34b7 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000010; // D (0x00000000000000000000000010000002) 
14'h212b : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000010; // D (0x00000000000000000000000020000002) 
14'h0a13 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000010; // D (0x00000000000000000000000040000002) 
14'h1f14 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000010; // D (0x00000000000000000000000080000002) 
14'h351a : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000010; // D (0x00000000000000000000000100000002) 
14'h2271 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000010; // D (0x00000000000000000000000200000002) 
14'h0ca7 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000010; // D (0x00000000000000000000000400000002) 
14'h127c : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000010; // D (0x00000000000000000000000800000002) 
14'h2fca : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000010; // D (0x00000000000000000000001000000002) 
14'h17d1 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000010; // D (0x00000000000000000000002000000002) 
14'h2490 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000010; // D (0x00000000000000000000004000000002) 
14'h0165 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000010; // D (0x00000000000000000000008000000002) 
14'h09f8 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000010; // D (0x00000000000000000000010000000002) 
14'h18c2 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000010; // D (0x00000000000000000000020000000002) 
14'h3ab6 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000010; // D (0x00000000000000000000040000000002) 
14'h3d29 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000010; // D (0x00000000000000000000080000000002) 
14'h3217 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000010; // D (0x00000000000000000000100000000002) 
14'h2c6b : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000010; // D (0x00000000000000000000200000000002) 
14'h1093 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000010; // D (0x00000000000000000000400000000002) 
14'h2a14 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000010; // D (0x00000000000000000000800000000002) 
14'h1c6d : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000010; // D (0x00000000000000000001000000000002) 
14'h33e8 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000010; // D (0x00000000000000000002000000000002) 
14'h2f95 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000010; // D (0x00000000000000000004000000000002) 
14'h176f : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000010; // D (0x00000000000000000008000000000002) 
14'h25ec : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000010; // D (0x00000000000000000010000000000002) 
14'h039d : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000010; // D (0x00000000000000000020000000000002) 
14'h0c08 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000010; // D (0x00000000000000000040000000000002) 
14'h1322 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000010; // D (0x00000000000000000080000000000002) 
14'h2d76 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000010; // D (0x00000000000000000100000000000002) 
14'h12a9 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000010; // D (0x00000000000000000200000000000002) 
14'h2e60 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000010; // D (0x00000000000000000400000000000002) 
14'h1485 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000010; // D (0x00000000000000000800000000000002) 
14'h2238 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000010; // D (0x00000000000000001000000000000002) 
14'h0c35 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000010; // D (0x00000000000000002000000000000002) 
14'h1358 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000010; // D (0x00000000000000004000000000000002) 
14'h2d82 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000010; // D (0x00000000000000008000000000000002) 
14'h1341 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000010; // D (0x00000000000000010000000000000002) 
14'h2db0 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000010; // D (0x00000000000000020000000000000002) 
14'h1325 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000010; // D (0x00000000000000040000000000000002) 
14'h2d78 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000010; // D (0x00000000000000080000000000000002) 
14'h12b5 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000010; // D (0x00000000000000100000000000000002) 
14'h2e58 : LOC =         127'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000010; // D (0x00000000000000200000000000000002) 
14'h14f5 : LOC =         127'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000010; // D (0x00000000000000400000000000000002) 
14'h22d8 : LOC =         127'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000010; // D (0x00000000000000800000000000000002) 
14'h0df5 : LOC =         127'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000010; // D (0x00000000000001000000000000000002) 
14'h10d8 : LOC =         127'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000010; // D (0x00000000000002000000000000000002) 
14'h2a82 : LOC =         127'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000010; // D (0x00000000000004000000000000000002) 
14'h1d41 : LOC =         127'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000010; // D (0x00000000000008000000000000000002) 
14'h31b0 : LOC =         127'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000010; // D (0x00000000000010000000000000000002) 
14'h2b25 : LOC =         127'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000010; // D (0x00000000000020000000000000000002) 
14'h1e0f : LOC =         127'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000010; // D (0x00000000000040000000000000000002) 
14'h372c : LOC =         127'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000010; // D (0x00000000000080000000000000000002) 
14'h261d : LOC =         127'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000010; // D (0x00000000000100000000000000000002) 
14'h047f : LOC =         127'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000010; // D (0x00000000000200000000000000000002) 
14'h03cc : LOC =         127'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000010; // D (0x00000000000400000000000000000002) 
14'h0caa : LOC =         127'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000010; // D (0x00000000000800000000000000000002) 
14'h1266 : LOC =         127'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000010; // D (0x00000000001000000000000000000002) 
14'h2ffe : LOC =         127'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000010; // D (0x00000000002000000000000000000002) 
14'h17b9 : LOC =         127'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000010; // D (0x00000000004000000000000000000002) 
14'h2440 : LOC =         127'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000010; // D (0x00000000008000000000000000000002) 
14'h00c5 : LOC =         127'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000010; // D (0x00000000010000000000000000000002) 
14'h0ab8 : LOC =         127'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000010; // D (0x00000000020000000000000000000002) 
14'h1e42 : LOC =         127'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010; // D (0x00000000040000000000000000000002) 
14'h37b6 : LOC =         127'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010; // D (0x00000000080000000000000000000002) 
14'h2729 : LOC =         127'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010; // D (0x00000000100000000000000000000002) 
14'h0617 : LOC =         127'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010; // D (0x00000000200000000000000000000002) 
14'h071c : LOC =         127'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010; // D (0x00000000400000000000000000000002) 
14'h050a : LOC =         127'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010; // D (0x00000000800000000000000000000002) 
14'h0126 : LOC =         127'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010; // D (0x00000001000000000000000000000002) 
14'h097e : LOC =         127'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010; // D (0x00000002000000000000000000000002) 
14'h19ce : LOC =         127'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010; // D (0x00000004000000000000000000000002) 
14'h38ae : LOC =         127'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010; // D (0x00000008000000000000000000000002) 
14'h3919 : LOC =         127'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010; // D (0x00000010000000000000000000000002) 
14'h3a77 : LOC =         127'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010; // D (0x00000020000000000000000000000002) 
14'h3cab : LOC =         127'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010; // D (0x00000040000000000000000000000002) 
14'h3113 : LOC =         127'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010; // D (0x00000080000000000000000000000002) 
14'h2a63 : LOC =         127'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010; // D (0x00000100000000000000000000000002) 
14'h1c83 : LOC =         127'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010; // D (0x00000200000000000000000000000002) 
14'h3234 : LOC =         127'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010; // D (0x00000400000000000000000000000002) 
14'h2c2d : LOC =         127'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010; // D (0x00000800000000000000000000000002) 
14'h101f : LOC =         127'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010; // D (0x00001000000000000000000000000002) 
14'h2b0c : LOC =         127'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010; // D (0x00002000000000000000000000000002) 
14'h1e5d : LOC =         127'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010; // D (0x00004000000000000000000000000002) 
14'h3788 : LOC =         127'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010; // D (0x00008000000000000000000000000002) 
14'h2755 : LOC =         127'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010; // D (0x00010000000000000000000000000002) 
14'h06ef : LOC =         127'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010; // D (0x00020000000000000000000000000002) 
14'h06ec : LOC =         127'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010; // D (0x00040000000000000000000000000002) 
14'h06ea : LOC =         127'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010; // D (0x00080000000000000000000000000002) 
14'h06e6 : LOC =         127'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010; // D (0x00100000000000000000000000000002) 
14'h06fe : LOC =         127'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010; // D (0x00200000000000000000000000000002) 
14'h06ce : LOC =         127'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010; // D (0x00400000000000000000000000000002) 
14'h06ae : LOC =         127'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010; // D (0x00800000000000000000000000000002) 
14'h066e : LOC =         127'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010; // D (0x01000000000000000000000000000002) 
14'h07ee : LOC =         127'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010; // D (0x02000000000000000000000000000002) 
14'h04ee : LOC =         127'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010; // D (0x04000000000000000000000000000002) 
14'h02ee : LOC =         127'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010; // D (0x08000000000000000000000000000002) 
14'h0eee : LOC =         127'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010; // D (0x10000000000000000000000000000002) 
14'h16ee : LOC =         127'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010; // D (0x20000000000000000000000000000002) 
14'h26ee : LOC =         127'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010; // D (0x40000000000000000000000000000002) 
14'h0ddc : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100; // S (0x00000000000000000000000000000004) 
14'h1664 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100; // D (0x0000000000000000000000000000000c) 
14'h3aac : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100; // D (0x00000000000000000000000000000014) 
14'h204b : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100; // D (0x00000000000000000000000000000024) 
14'h1585 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000100; // D (0x00000000000000000000000000000044) 
14'h3d6e : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000100; // D (0x00000000000000000000000000000084) 
14'h2fcf : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000100; // D (0x00000000000000000000000000000104) 
14'h0a8d : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000100; // D (0x00000000000000000000000000000204) 
14'h037e : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000100; // D (0x00000000000000000000000000000404) 
14'h1098 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000100; // D (0x00000000000000000000000000000804) 
14'h3754 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000100; // D (0x00000000000000000000000000001004) 
14'h3bbb : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000100; // D (0x00000000000000000000000000002004) 
14'h2265 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000100; // D (0x00000000000000000000000000004004) 
14'h11d9 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000100; // D (0x00000000000000000000000000008004) 
14'h35d6 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000100; // D (0x00000000000000000000000000010004) 
14'h3ebf : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000100; // D (0x00000000000000000000000000020004) 
14'h286d : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000100; // D (0x00000000000000000000000000040004) 
14'h05c9 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000100; // D (0x00000000000000000000000000080004) 
14'h1df6 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000100; // D (0x00000000000000000000000000100004) 
14'h2d88 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000100; // D (0x00000000000000000000000000200004) 
14'h0e03 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000100; // D (0x00000000000000000000000000400004) 
14'h0a62 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000100; // D (0x00000000000000000000000000800004) 
14'h02a0 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000100; // D (0x00000000000000000000000001000004) 
14'h1324 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000100; // D (0x00000000000000000000000002000004) 
14'h302c : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000100; // D (0x00000000000000000000000004000004) 
14'h354b : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000100; // D (0x00000000000000000000000008000004) 
14'h3f85 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000100; // D (0x00000000000000000000000010000004) 
14'h2a19 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000100; // D (0x00000000000000000000000020000004) 
14'h0121 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000100; // D (0x00000000000000000000000040000004) 
14'h1426 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000100; // D (0x00000000000000000000000080000004) 
14'h3e28 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000100; // D (0x00000000000000000000000100000004) 
14'h2943 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000100; // D (0x00000000000000000000000200000004) 
14'h0795 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000100; // D (0x00000000000000000000000400000004) 
14'h194e : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000100; // D (0x00000000000000000000000800000004) 
14'h24f8 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000100; // D (0x00000000000000000000001000000004) 
14'h1ce3 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000100; // D (0x00000000000000000000002000000004) 
14'h2fa2 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000100; // D (0x00000000000000000000004000000004) 
14'h0a57 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000100; // D (0x00000000000000000000008000000004) 
14'h02ca : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000100; // D (0x00000000000000000000010000000004) 
14'h13f0 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000100; // D (0x00000000000000000000020000000004) 
14'h3184 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000100; // D (0x00000000000000000000040000000004) 
14'h361b : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000100; // D (0x00000000000000000000080000000004) 
14'h3925 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000100; // D (0x00000000000000000000100000000004) 
14'h2759 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000100; // D (0x00000000000000000000200000000004) 
14'h1ba1 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000100; // D (0x00000000000000000000400000000004) 
14'h2126 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000100; // D (0x00000000000000000000800000000004) 
14'h175f : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000100; // D (0x00000000000000000001000000000004) 
14'h38da : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000100; // D (0x00000000000000000002000000000004) 
14'h24a7 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000100; // D (0x00000000000000000004000000000004) 
14'h1c5d : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000100; // D (0x00000000000000000008000000000004) 
14'h2ede : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000100; // D (0x00000000000000000010000000000004) 
14'h08af : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000100; // D (0x00000000000000000020000000000004) 
14'h073a : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000100; // D (0x00000000000000000040000000000004) 
14'h1810 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000100; // D (0x00000000000000000080000000000004) 
14'h2644 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000100; // D (0x00000000000000000100000000000004) 
14'h199b : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000100; // D (0x00000000000000000200000000000004) 
14'h2552 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000100; // D (0x00000000000000000400000000000004) 
14'h1fb7 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000100; // D (0x00000000000000000800000000000004) 
14'h290a : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000100; // D (0x00000000000000001000000000000004) 
14'h0707 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000100; // D (0x00000000000000002000000000000004) 
14'h186a : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000100; // D (0x00000000000000004000000000000004) 
14'h26b0 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000100; // D (0x00000000000000008000000000000004) 
14'h1873 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000100; // D (0x00000000000000010000000000000004) 
14'h2682 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000100; // D (0x00000000000000020000000000000004) 
14'h1817 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000100; // D (0x00000000000000040000000000000004) 
14'h264a : LOC =         127'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000100; // D (0x00000000000000080000000000000004) 
14'h1987 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000100; // D (0x00000000000000100000000000000004) 
14'h256a : LOC =         127'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000100; // D (0x00000000000000200000000000000004) 
14'h1fc7 : LOC =         127'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000100; // D (0x00000000000000400000000000000004) 
14'h29ea : LOC =         127'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000100; // D (0x00000000000000800000000000000004) 
14'h06c7 : LOC =         127'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000100; // D (0x00000000000001000000000000000004) 
14'h1bea : LOC =         127'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000100; // D (0x00000000000002000000000000000004) 
14'h21b0 : LOC =         127'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000100; // D (0x00000000000004000000000000000004) 
14'h1673 : LOC =         127'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000100; // D (0x00000000000008000000000000000004) 
14'h3a82 : LOC =         127'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000100; // D (0x00000000000010000000000000000004) 
14'h2017 : LOC =         127'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000100; // D (0x00000000000020000000000000000004) 
14'h153d : LOC =         127'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000100; // D (0x00000000000040000000000000000004) 
14'h3c1e : LOC =         127'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000100; // D (0x00000000000080000000000000000004) 
14'h2d2f : LOC =         127'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000100; // D (0x00000000000100000000000000000004) 
14'h0f4d : LOC =         127'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000100; // D (0x00000000000200000000000000000004) 
14'h08fe : LOC =         127'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000100; // D (0x00000000000400000000000000000004) 
14'h0798 : LOC =         127'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000100; // D (0x00000000000800000000000000000004) 
14'h1954 : LOC =         127'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000100; // D (0x00000000001000000000000000000004) 
14'h24cc : LOC =         127'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100; // D (0x00000000002000000000000000000004) 
14'h1c8b : LOC =         127'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000100; // D (0x00000000004000000000000000000004) 
14'h2f72 : LOC =         127'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000100; // D (0x00000000008000000000000000000004) 
14'h0bf7 : LOC =         127'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000100; // D (0x00000000010000000000000000000004) 
14'h018a : LOC =         127'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000100; // D (0x00000000020000000000000000000004) 
14'h1570 : LOC =         127'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100; // D (0x00000000040000000000000000000004) 
14'h3c84 : LOC =         127'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100; // D (0x00000000080000000000000000000004) 
14'h2c1b : LOC =         127'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100; // D (0x00000000100000000000000000000004) 
14'h0d25 : LOC =         127'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100; // D (0x00000000200000000000000000000004) 
14'h0c2e : LOC =         127'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100; // D (0x00000000400000000000000000000004) 
14'h0e38 : LOC =         127'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100; // D (0x00000000800000000000000000000004) 
14'h0a14 : LOC =         127'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100; // D (0x00000001000000000000000000000004) 
14'h024c : LOC =         127'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100; // D (0x00000002000000000000000000000004) 
14'h12fc : LOC =         127'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100; // D (0x00000004000000000000000000000004) 
14'h339c : LOC =         127'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100; // D (0x00000008000000000000000000000004) 
14'h322b : LOC =         127'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100; // D (0x00000010000000000000000000000004) 
14'h3145 : LOC =         127'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100; // D (0x00000020000000000000000000000004) 
14'h3799 : LOC =         127'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100; // D (0x00000040000000000000000000000004) 
14'h3a21 : LOC =         127'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100; // D (0x00000080000000000000000000000004) 
14'h2151 : LOC =         127'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100; // D (0x00000100000000000000000000000004) 
14'h17b1 : LOC =         127'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100; // D (0x00000200000000000000000000000004) 
14'h3906 : LOC =         127'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100; // D (0x00000400000000000000000000000004) 
14'h271f : LOC =         127'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100; // D (0x00000800000000000000000000000004) 
14'h1b2d : LOC =         127'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100; // D (0x00001000000000000000000000000004) 
14'h203e : LOC =         127'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100; // D (0x00002000000000000000000000000004) 
14'h156f : LOC =         127'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100; // D (0x00004000000000000000000000000004) 
14'h3cba : LOC =         127'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100; // D (0x00008000000000000000000000000004) 
14'h2c67 : LOC =         127'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100; // D (0x00010000000000000000000000000004) 
14'h0ddd : LOC =         127'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100; // D (0x00020000000000000000000000000004) 
14'h0dde : LOC =         127'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100; // D (0x00040000000000000000000000000004) 
14'h0dd8 : LOC =         127'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100; // D (0x00080000000000000000000000000004) 
14'h0dd4 : LOC =         127'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100; // D (0x00100000000000000000000000000004) 
14'h0dcc : LOC =         127'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100; // D (0x00200000000000000000000000000004) 
14'h0dfc : LOC =         127'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100; // D (0x00400000000000000000000000000004) 
14'h0d9c : LOC =         127'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100; // D (0x00800000000000000000000000000004) 
14'h0d5c : LOC =         127'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100; // D (0x01000000000000000000000000000004) 
14'h0cdc : LOC =         127'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100; // D (0x02000000000000000000000000000004) 
14'h0fdc : LOC =         127'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100; // D (0x04000000000000000000000000000004) 
14'h09dc : LOC =         127'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100; // D (0x08000000000000000000000000000004) 
14'h05dc : LOC =         127'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100; // D (0x10000000000000000000000000000004) 
14'h1ddc : LOC =         127'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100; // D (0x20000000000000000000000000000004) 
14'h2ddc : LOC =         127'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100; // D (0x40000000000000000000000000000004) 
14'h1bb8 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000; // S (0x00000000000000000000000000000008) 
14'h2cc8 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000; // D (0x00000000000000000000000000000018) 
14'h362f : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000; // D (0x00000000000000000000000000000028) 
14'h03e1 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000; // D (0x00000000000000000000000000000048) 
14'h2b0a : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000; // D (0x00000000000000000000000000000088) 
14'h39ab : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100001000; // D (0x00000000000000000000000000000108) 
14'h1ce9 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000001000; // D (0x00000000000000000000000000000208) 
14'h151a : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000001000; // D (0x00000000000000000000000000000408) 
14'h06fc : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000001000; // D (0x00000000000000000000000000000808) 
14'h2130 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000001000; // D (0x00000000000000000000000000001008) 
14'h2ddf : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000001000; // D (0x00000000000000000000000000002008) 
14'h3401 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000001000; // D (0x00000000000000000000000000004008) 
14'h07bd : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000001000; // D (0x00000000000000000000000000008008) 
14'h23b2 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000001000; // D (0x00000000000000000000000000010008) 
14'h28db : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000001000; // D (0x00000000000000000000000000020008) 
14'h3e09 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000001000; // D (0x00000000000000000000000000040008) 
14'h13ad : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001000; // D (0x00000000000000000000000000080008) 
14'h0b92 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000001000; // D (0x00000000000000000000000000100008) 
14'h3bec : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000001000; // D (0x00000000000000000000000000200008) 
14'h1867 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000001000; // D (0x00000000000000000000000000400008) 
14'h1c06 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000001000; // D (0x00000000000000000000000000800008) 
14'h14c4 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000001000; // D (0x00000000000000000000000001000008) 
14'h0540 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000001000; // D (0x00000000000000000000000002000008) 
14'h2648 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000001000; // D (0x00000000000000000000000004000008) 
14'h232f : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000001000; // D (0x00000000000000000000000008000008) 
14'h29e1 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000001000; // D (0x00000000000000000000000010000008) 
14'h3c7d : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000001000; // D (0x00000000000000000000000020000008) 
14'h1745 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000001000; // D (0x00000000000000000000000040000008) 
14'h0242 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000001000; // D (0x00000000000000000000000080000008) 
14'h284c : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000001000; // D (0x00000000000000000000000100000008) 
14'h3f27 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000001000; // D (0x00000000000000000000000200000008) 
14'h11f1 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000001000; // D (0x00000000000000000000000400000008) 
14'h0f2a : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000001000; // D (0x00000000000000000000000800000008) 
14'h329c : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000001000; // D (0x00000000000000000000001000000008) 
14'h0a87 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000001000; // D (0x00000000000000000000002000000008) 
14'h39c6 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000001000; // D (0x00000000000000000000004000000008) 
14'h1c33 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000001000; // D (0x00000000000000000000008000000008) 
14'h14ae : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000001000; // D (0x00000000000000000000010000000008) 
14'h0594 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000001000; // D (0x00000000000000000000020000000008) 
14'h27e0 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000001000; // D (0x00000000000000000000040000000008) 
14'h207f : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000001000; // D (0x00000000000000000000080000000008) 
14'h2f41 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000001000; // D (0x00000000000000000000100000000008) 
14'h313d : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000001000; // D (0x00000000000000000000200000000008) 
14'h0dc5 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000001000; // D (0x00000000000000000000400000000008) 
14'h3742 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000001000; // D (0x00000000000000000000800000000008) 
14'h013b : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000001000; // D (0x00000000000000000001000000000008) 
14'h2ebe : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000001000; // D (0x00000000000000000002000000000008) 
14'h32c3 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000001000; // D (0x00000000000000000004000000000008) 
14'h0a39 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000001000; // D (0x00000000000000000008000000000008) 
14'h38ba : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000001000; // D (0x00000000000000000010000000000008) 
14'h1ecb : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000001000; // D (0x00000000000000000020000000000008) 
14'h115e : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000001000; // D (0x00000000000000000040000000000008) 
14'h0e74 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000001000; // D (0x00000000000000000080000000000008) 
14'h3020 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000001000; // D (0x00000000000000000100000000000008) 
14'h0fff : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000001000; // D (0x00000000000000000200000000000008) 
14'h3336 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000001000; // D (0x00000000000000000400000000000008) 
14'h09d3 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000001000; // D (0x00000000000000000800000000000008) 
14'h3f6e : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000001000; // D (0x00000000000000001000000000000008) 
14'h1163 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000001000; // D (0x00000000000000002000000000000008) 
14'h0e0e : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000001000; // D (0x00000000000000004000000000000008) 
14'h30d4 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000001000; // D (0x00000000000000008000000000000008) 
14'h0e17 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000001000; // D (0x00000000000000010000000000000008) 
14'h30e6 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000001000; // D (0x00000000000000020000000000000008) 
14'h0e73 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000001000; // D (0x00000000000000040000000000000008) 
14'h302e : LOC =         127'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000001000; // D (0x00000000000000080000000000000008) 
14'h0fe3 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000001000; // D (0x00000000000000100000000000000008) 
14'h330e : LOC =         127'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000001000; // D (0x00000000000000200000000000000008) 
14'h09a3 : LOC =         127'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000001000; // D (0x00000000000000400000000000000008) 
14'h3f8e : LOC =         127'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000001000; // D (0x00000000000000800000000000000008) 
14'h10a3 : LOC =         127'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000001000; // D (0x00000000000001000000000000000008) 
14'h0d8e : LOC =         127'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000001000; // D (0x00000000000002000000000000000008) 
14'h37d4 : LOC =         127'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000001000; // D (0x00000000000004000000000000000008) 
14'h0017 : LOC =         127'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000001000; // D (0x00000000000008000000000000000008) 
14'h2ce6 : LOC =         127'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000001000; // D (0x00000000000010000000000000000008) 
14'h3673 : LOC =         127'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000001000; // D (0x00000000000020000000000000000008) 
14'h0359 : LOC =         127'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000001000; // D (0x00000000000040000000000000000008) 
14'h2a7a : LOC =         127'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000001000; // D (0x00000000000080000000000000000008) 
14'h3b4b : LOC =         127'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000001000; // D (0x00000000000100000000000000000008) 
14'h1929 : LOC =         127'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000001000; // D (0x00000000000200000000000000000008) 
14'h1e9a : LOC =         127'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000001000; // D (0x00000000000400000000000000000008) 
14'h11fc : LOC =         127'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000001000; // D (0x00000000000800000000000000000008) 
14'h0f30 : LOC =         127'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000001000; // D (0x00000000001000000000000000000008) 
14'h32a8 : LOC =         127'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000001000; // D (0x00000000002000000000000000000008) 
14'h0aef : LOC =         127'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000001000; // D (0x00000000004000000000000000000008) 
14'h3916 : LOC =         127'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000001000; // D (0x00000000008000000000000000000008) 
14'h1d93 : LOC =         127'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000001000; // D (0x00000000010000000000000000000008) 
14'h17ee : LOC =         127'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000001000; // D (0x00000000020000000000000000000008) 
14'h0314 : LOC =         127'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000; // D (0x00000000040000000000000000000008) 
14'h2ae0 : LOC =         127'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000; // D (0x00000000080000000000000000000008) 
14'h3a7f : LOC =         127'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000; // D (0x00000000100000000000000000000008) 
14'h1b41 : LOC =         127'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000; // D (0x00000000200000000000000000000008) 
14'h1a4a : LOC =         127'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000; // D (0x00000000400000000000000000000008) 
14'h185c : LOC =         127'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000; // D (0x00000000800000000000000000000008) 
14'h1c70 : LOC =         127'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000; // D (0x00000001000000000000000000000008) 
14'h1428 : LOC =         127'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000; // D (0x00000002000000000000000000000008) 
14'h0498 : LOC =         127'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000; // D (0x00000004000000000000000000000008) 
14'h25f8 : LOC =         127'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000; // D (0x00000008000000000000000000000008) 
14'h244f : LOC =         127'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000; // D (0x00000010000000000000000000000008) 
14'h2721 : LOC =         127'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000; // D (0x00000020000000000000000000000008) 
14'h21fd : LOC =         127'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000; // D (0x00000040000000000000000000000008) 
14'h2c45 : LOC =         127'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000; // D (0x00000080000000000000000000000008) 
14'h3735 : LOC =         127'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000; // D (0x00000100000000000000000000000008) 
14'h01d5 : LOC =         127'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000; // D (0x00000200000000000000000000000008) 
14'h2f62 : LOC =         127'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000; // D (0x00000400000000000000000000000008) 
14'h317b : LOC =         127'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000; // D (0x00000800000000000000000000000008) 
14'h0d49 : LOC =         127'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000; // D (0x00001000000000000000000000000008) 
14'h365a : LOC =         127'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000; // D (0x00002000000000000000000000000008) 
14'h030b : LOC =         127'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000; // D (0x00004000000000000000000000000008) 
14'h2ade : LOC =         127'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000; // D (0x00008000000000000000000000000008) 
14'h3a03 : LOC =         127'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000; // D (0x00010000000000000000000000000008) 
14'h1bb9 : LOC =         127'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000; // D (0x00020000000000000000000000000008) 
14'h1bba : LOC =         127'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000; // D (0x00040000000000000000000000000008) 
14'h1bbc : LOC =         127'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000; // D (0x00080000000000000000000000000008) 
14'h1bb0 : LOC =         127'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000; // D (0x00100000000000000000000000000008) 
14'h1ba8 : LOC =         127'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000; // D (0x00200000000000000000000000000008) 
14'h1b98 : LOC =         127'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000; // D (0x00400000000000000000000000000008) 
14'h1bf8 : LOC =         127'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000; // D (0x00800000000000000000000000000008) 
14'h1b38 : LOC =         127'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000; // D (0x01000000000000000000000000000008) 
14'h1ab8 : LOC =         127'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000; // D (0x02000000000000000000000000000008) 
14'h19b8 : LOC =         127'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000; // D (0x04000000000000000000000000000008) 
14'h1fb8 : LOC =         127'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000; // D (0x08000000000000000000000000000008) 
14'h13b8 : LOC =         127'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000; // D (0x10000000000000000000000000000008) 
14'h0bb8 : LOC =         127'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000; // D (0x20000000000000000000000000000008) 
14'h3bb8 : LOC =         127'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000; // D (0x40000000000000000000000000000008) 
14'h3770 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000; // S (0x00000000000000000000000000000010) 
14'h1ae7 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000; // D (0x00000000000000000000000000000030) 
14'h2f29 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000; // D (0x00000000000000000000000000000050) 
14'h07c2 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000; // D (0x00000000000000000000000000000090) 
14'h1563 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010000; // D (0x00000000000000000000000000000110) 
14'h3021 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000010000; // D (0x00000000000000000000000000000210) 
14'h39d2 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000010000; // D (0x00000000000000000000000000000410) 
14'h2a34 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000010000; // D (0x00000000000000000000000000000810) 
14'h0df8 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000010000; // D (0x00000000000000000000000000001010) 
14'h0117 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000010000; // D (0x00000000000000000000000000002010) 
14'h18c9 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000010000; // D (0x00000000000000000000000000004010) 
14'h2b75 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000010000; // D (0x00000000000000000000000000008010) 
14'h0f7a : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000010000; // D (0x00000000000000000000000000010010) 
14'h0413 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000010000; // D (0x00000000000000000000000000020010) 
14'h12c1 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000010000; // D (0x00000000000000000000000000040010) 
14'h3f65 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000010000; // D (0x00000000000000000000000000080010) 
14'h275a : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000010000; // D (0x00000000000000000000000000100010) 
14'h1724 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000010000; // D (0x00000000000000000000000000200010) 
14'h34af : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000010000; // D (0x00000000000000000000000000400010) 
14'h30ce : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000010000; // D (0x00000000000000000000000000800010) 
14'h380c : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000010000; // D (0x00000000000000000000000001000010) 
14'h2988 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000010000; // D (0x00000000000000000000000002000010) 
14'h0a80 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000010000; // D (0x00000000000000000000000004000010) 
14'h0fe7 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000010000; // D (0x00000000000000000000000008000010) 
14'h0529 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000010000; // D (0x00000000000000000000000010000010) 
14'h10b5 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000010000; // D (0x00000000000000000000000020000010) 
14'h3b8d : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000010000; // D (0x00000000000000000000000040000010) 
14'h2e8a : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000010000; // D (0x00000000000000000000000080000010) 
14'h0484 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000010000; // D (0x00000000000000000000000100000010) 
14'h13ef : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000010000; // D (0x00000000000000000000000200000010) 
14'h3d39 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000010000; // D (0x00000000000000000000000400000010) 
14'h23e2 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000010000; // D (0x00000000000000000000000800000010) 
14'h1e54 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000010000; // D (0x00000000000000000000001000000010) 
14'h264f : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000010000; // D (0x00000000000000000000002000000010) 
14'h150e : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000010000; // D (0x00000000000000000000004000000010) 
14'h30fb : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000010000; // D (0x00000000000000000000008000000010) 
14'h3866 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000010000; // D (0x00000000000000000000010000000010) 
14'h295c : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000010000; // D (0x00000000000000000000020000000010) 
14'h0b28 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000010000; // D (0x00000000000000000000040000000010) 
14'h0cb7 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000010000; // D (0x00000000000000000000080000000010) 
14'h0389 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000010000; // D (0x00000000000000000000100000000010) 
14'h1df5 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000010000; // D (0x00000000000000000000200000000010) 
14'h210d : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000010000; // D (0x00000000000000000000400000000010) 
14'h1b8a : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000010000; // D (0x00000000000000000000800000000010) 
14'h2df3 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000010000; // D (0x00000000000000000001000000000010) 
14'h0276 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000010000; // D (0x00000000000000000002000000000010) 
14'h1e0b : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000010000; // D (0x00000000000000000004000000000010) 
14'h26f1 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000010000; // D (0x00000000000000000008000000000010) 
14'h1472 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000010000; // D (0x00000000000000000010000000000010) 
14'h3203 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000010000; // D (0x00000000000000000020000000000010) 
14'h3d96 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000010000; // D (0x00000000000000000040000000000010) 
14'h22bc : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000010000; // D (0x00000000000000000080000000000010) 
14'h1ce8 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000010000; // D (0x00000000000000000100000000000010) 
14'h2337 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000010000; // D (0x00000000000000000200000000000010) 
14'h1ffe : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000010000; // D (0x00000000000000000400000000000010) 
14'h251b : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000010000; // D (0x00000000000000000800000000000010) 
14'h13a6 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000010000; // D (0x00000000000000001000000000000010) 
14'h3dab : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000010000; // D (0x00000000000000002000000000000010) 
14'h22c6 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000010000; // D (0x00000000000000004000000000000010) 
14'h1c1c : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000010000; // D (0x00000000000000008000000000000010) 
14'h22df : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000010000; // D (0x00000000000000010000000000000010) 
14'h1c2e : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000010000; // D (0x00000000000000020000000000000010) 
14'h22bb : LOC =         127'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000010000; // D (0x00000000000000040000000000000010) 
14'h1ce6 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000010000; // D (0x00000000000000080000000000000010) 
14'h232b : LOC =         127'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000010000; // D (0x00000000000000100000000000000010) 
14'h1fc6 : LOC =         127'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000010000; // D (0x00000000000000200000000000000010) 
14'h256b : LOC =         127'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000010000; // D (0x00000000000000400000000000000010) 
14'h1346 : LOC =         127'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000010000; // D (0x00000000000000800000000000000010) 
14'h3c6b : LOC =         127'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000010000; // D (0x00000000000001000000000000000010) 
14'h2146 : LOC =         127'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000010000; // D (0x00000000000002000000000000000010) 
14'h1b1c : LOC =         127'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000010000; // D (0x00000000000004000000000000000010) 
14'h2cdf : LOC =         127'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000010000; // D (0x00000000000008000000000000000010) 
14'h002e : LOC =         127'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000010000; // D (0x00000000000010000000000000000010) 
14'h1abb : LOC =         127'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000010000; // D (0x00000000000020000000000000000010) 
14'h2f91 : LOC =         127'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000010000; // D (0x00000000000040000000000000000010) 
14'h06b2 : LOC =         127'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000010000; // D (0x00000000000080000000000000000010) 
14'h1783 : LOC =         127'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000010000; // D (0x00000000000100000000000000000010) 
14'h35e1 : LOC =         127'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000010000; // D (0x00000000000200000000000000000010) 
14'h3252 : LOC =         127'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000010000; // D (0x00000000000400000000000000000010) 
14'h3d34 : LOC =         127'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000010000; // D (0x00000000000800000000000000000010) 
14'h23f8 : LOC =         127'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000010000; // D (0x00000000001000000000000000000010) 
14'h1e60 : LOC =         127'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000010000; // D (0x00000000002000000000000000000010) 
14'h2627 : LOC =         127'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000010000; // D (0x00000000004000000000000000000010) 
14'h15de : LOC =         127'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000010000; // D (0x00000000008000000000000000000010) 
14'h315b : LOC =         127'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000010000; // D (0x00000000010000000000000000000010) 
14'h3b26 : LOC =         127'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000010000; // D (0x00000000020000000000000000000010) 
14'h2fdc : LOC =         127'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000; // D (0x00000000040000000000000000000010) 
14'h0628 : LOC =         127'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000; // D (0x00000000080000000000000000000010) 
14'h16b7 : LOC =         127'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000; // D (0x00000000100000000000000000000010) 
14'h3789 : LOC =         127'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000; // D (0x00000000200000000000000000000010) 
14'h3682 : LOC =         127'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000; // D (0x00000000400000000000000000000010) 
14'h3494 : LOC =         127'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000; // D (0x00000000800000000000000000000010) 
14'h30b8 : LOC =         127'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000; // D (0x00000001000000000000000000000010) 
14'h38e0 : LOC =         127'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000; // D (0x00000002000000000000000000000010) 
14'h2850 : LOC =         127'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000; // D (0x00000004000000000000000000000010) 
14'h0930 : LOC =         127'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000; // D (0x00000008000000000000000000000010) 
14'h0887 : LOC =         127'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000; // D (0x00000010000000000000000000000010) 
14'h0be9 : LOC =         127'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000; // D (0x00000020000000000000000000000010) 
14'h0d35 : LOC =         127'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000; // D (0x00000040000000000000000000000010) 
14'h008d : LOC =         127'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000; // D (0x00000080000000000000000000000010) 
14'h1bfd : LOC =         127'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000; // D (0x00000100000000000000000000000010) 
14'h2d1d : LOC =         127'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000; // D (0x00000200000000000000000000000010) 
14'h03aa : LOC =         127'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000; // D (0x00000400000000000000000000000010) 
14'h1db3 : LOC =         127'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000; // D (0x00000800000000000000000000000010) 
14'h2181 : LOC =         127'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000; // D (0x00001000000000000000000000000010) 
14'h1a92 : LOC =         127'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000; // D (0x00002000000000000000000000000010) 
14'h2fc3 : LOC =         127'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000; // D (0x00004000000000000000000000000010) 
14'h0616 : LOC =         127'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000; // D (0x00008000000000000000000000000010) 
14'h16cb : LOC =         127'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000; // D (0x00010000000000000000000000000010) 
14'h3771 : LOC =         127'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000; // D (0x00020000000000000000000000000010) 
14'h3772 : LOC =         127'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000; // D (0x00040000000000000000000000000010) 
14'h3774 : LOC =         127'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000; // D (0x00080000000000000000000000000010) 
14'h3778 : LOC =         127'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000; // D (0x00100000000000000000000000000010) 
14'h3760 : LOC =         127'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000; // D (0x00200000000000000000000000000010) 
14'h3750 : LOC =         127'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000; // D (0x00400000000000000000000000000010) 
14'h3730 : LOC =         127'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000; // D (0x00800000000000000000000000000010) 
14'h37f0 : LOC =         127'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000; // D (0x01000000000000000000000000000010) 
14'h3670 : LOC =         127'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000; // D (0x02000000000000000000000000000010) 
14'h3570 : LOC =         127'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000; // D (0x04000000000000000000000000000010) 
14'h3370 : LOC =         127'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000; // D (0x08000000000000000000000000000010) 
14'h3f70 : LOC =         127'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000; // D (0x10000000000000000000000000000010) 
14'h2770 : LOC =         127'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000; // D (0x20000000000000000000000000000010) 
14'h1770 : LOC =         127'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000; // D (0x40000000000000000000000000000010) 
14'h2d97 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000; // S (0x00000000000000000000000000000020) 
14'h35ce : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000; // D (0x00000000000000000000000000000060) 
14'h1d25 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000; // D (0x000000000000000000000000000000a0) 
14'h0f84 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000; // D (0x00000000000000000000000000000120) 
14'h2ac6 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000100000; // D (0x00000000000000000000000000000220) 
14'h2335 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000100000; // D (0x00000000000000000000000000000420) 
14'h30d3 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000100000; // D (0x00000000000000000000000000000820) 
14'h171f : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000100000; // D (0x00000000000000000000000000001020) 
14'h1bf0 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000100000; // D (0x00000000000000000000000000002020) 
14'h022e : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000100000; // D (0x00000000000000000000000000004020) 
14'h3192 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000100000; // D (0x00000000000000000000000000008020) 
14'h159d : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000100000; // D (0x00000000000000000000000000010020) 
14'h1ef4 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000100000; // D (0x00000000000000000000000000020020) 
14'h0826 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000100000; // D (0x00000000000000000000000000040020) 
14'h2582 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000100000; // D (0x00000000000000000000000000080020) 
14'h3dbd : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000100000; // D (0x00000000000000000000000000100020) 
14'h0dc3 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000100000; // D (0x00000000000000000000000000200020) 
14'h2e48 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000100000; // D (0x00000000000000000000000000400020) 
14'h2a29 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000100000; // D (0x00000000000000000000000000800020) 
14'h22eb : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000100000; // D (0x00000000000000000000000001000020) 
14'h336f : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000100000; // D (0x00000000000000000000000002000020) 
14'h1067 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000100000; // D (0x00000000000000000000000004000020) 
14'h1500 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000100000; // D (0x00000000000000000000000008000020) 
14'h1fce : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000100000; // D (0x00000000000000000000000010000020) 
14'h0a52 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000100000; // D (0x00000000000000000000000020000020) 
14'h216a : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000100000; // D (0x00000000000000000000000040000020) 
14'h346d : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000100000; // D (0x00000000000000000000000080000020) 
14'h1e63 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000100000; // D (0x00000000000000000000000100000020) 
14'h0908 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000100000; // D (0x00000000000000000000000200000020) 
14'h27de : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000100000; // D (0x00000000000000000000000400000020) 
14'h3905 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000100000; // D (0x00000000000000000000000800000020) 
14'h04b3 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000100000; // D (0x00000000000000000000001000000020) 
14'h3ca8 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000100000; // D (0x00000000000000000000002000000020) 
14'h0fe9 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000100000; // D (0x00000000000000000000004000000020) 
14'h2a1c : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000100000; // D (0x00000000000000000000008000000020) 
14'h2281 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000100000; // D (0x00000000000000000000010000000020) 
14'h33bb : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000100000; // D (0x00000000000000000000020000000020) 
14'h11cf : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000100000; // D (0x00000000000000000000040000000020) 
14'h1650 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000100000; // D (0x00000000000000000000080000000020) 
14'h196e : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000100000; // D (0x00000000000000000000100000000020) 
14'h0712 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000100000; // D (0x00000000000000000000200000000020) 
14'h3bea : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000100000; // D (0x00000000000000000000400000000020) 
14'h016d : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000100000; // D (0x00000000000000000000800000000020) 
14'h3714 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000100000; // D (0x00000000000000000001000000000020) 
14'h1891 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000100000; // D (0x00000000000000000002000000000020) 
14'h04ec : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000100000; // D (0x00000000000000000004000000000020) 
14'h3c16 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000100000; // D (0x00000000000000000008000000000020) 
14'h0e95 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000100000; // D (0x00000000000000000010000000000020) 
14'h28e4 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000100000; // D (0x00000000000000000020000000000020) 
14'h2771 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000100000; // D (0x00000000000000000040000000000020) 
14'h385b : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000100000; // D (0x00000000000000000080000000000020) 
14'h060f : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000100000; // D (0x00000000000000000100000000000020) 
14'h39d0 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000100000; // D (0x00000000000000000200000000000020) 
14'h0519 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000100000; // D (0x00000000000000000400000000000020) 
14'h3ffc : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000100000; // D (0x00000000000000000800000000000020) 
14'h0941 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000100000; // D (0x00000000000000001000000000000020) 
14'h274c : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000100000; // D (0x00000000000000002000000000000020) 
14'h3821 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000100000; // D (0x00000000000000004000000000000020) 
14'h06fb : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000100000; // D (0x00000000000000008000000000000020) 
14'h3838 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000100000; // D (0x00000000000000010000000000000020) 
14'h06c9 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000100000; // D (0x00000000000000020000000000000020) 
14'h385c : LOC =         127'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000100000; // D (0x00000000000000040000000000000020) 
14'h0601 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000100000; // D (0x00000000000000080000000000000020) 
14'h39cc : LOC =         127'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000100000; // D (0x00000000000000100000000000000020) 
14'h0521 : LOC =         127'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000100000; // D (0x00000000000000200000000000000020) 
14'h3f8c : LOC =         127'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000100000; // D (0x00000000000000400000000000000020) 
14'h09a1 : LOC =         127'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000100000; // D (0x00000000000000800000000000000020) 
14'h268c : LOC =         127'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000100000; // D (0x00000000000001000000000000000020) 
14'h3ba1 : LOC =         127'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000100000; // D (0x00000000000002000000000000000020) 
14'h01fb : LOC =         127'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000100000; // D (0x00000000000004000000000000000020) 
14'h3638 : LOC =         127'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000100000; // D (0x00000000000008000000000000000020) 
14'h1ac9 : LOC =         127'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000100000; // D (0x00000000000010000000000000000020) 
14'h005c : LOC =         127'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000100000; // D (0x00000000000020000000000000000020) 
14'h3576 : LOC =         127'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000100000; // D (0x00000000000040000000000000000020) 
14'h1c55 : LOC =         127'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000100000; // D (0x00000000000080000000000000000020) 
14'h0d64 : LOC =         127'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000100000; // D (0x00000000000100000000000000000020) 
14'h2f06 : LOC =         127'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000100000; // D (0x00000000000200000000000000000020) 
14'h28b5 : LOC =         127'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000100000; // D (0x00000000000400000000000000000020) 
14'h27d3 : LOC =         127'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000100000; // D (0x00000000000800000000000000000020) 
14'h391f : LOC =         127'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000100000; // D (0x00000000001000000000000000000020) 
14'h0487 : LOC =         127'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000100000; // D (0x00000000002000000000000000000020) 
14'h3cc0 : LOC =         127'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000100000; // D (0x00000000004000000000000000000020) 
14'h0f39 : LOC =         127'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000100000; // D (0x00000000008000000000000000000020) 
14'h2bbc : LOC =         127'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000; // D (0x00000000010000000000000000000020) 
14'h21c1 : LOC =         127'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000100000; // D (0x00000000020000000000000000000020) 
14'h353b : LOC =         127'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000; // D (0x00000000040000000000000000000020) 
14'h1ccf : LOC =         127'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000; // D (0x00000000080000000000000000000020) 
14'h0c50 : LOC =         127'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000; // D (0x00000000100000000000000000000020) 
14'h2d6e : LOC =         127'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000; // D (0x00000000200000000000000000000020) 
14'h2c65 : LOC =         127'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000; // D (0x00000000400000000000000000000020) 
14'h2e73 : LOC =         127'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000; // D (0x00000000800000000000000000000020) 
14'h2a5f : LOC =         127'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000; // D (0x00000001000000000000000000000020) 
14'h2207 : LOC =         127'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000; // D (0x00000002000000000000000000000020) 
14'h32b7 : LOC =         127'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000; // D (0x00000004000000000000000000000020) 
14'h13d7 : LOC =         127'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000; // D (0x00000008000000000000000000000020) 
14'h1260 : LOC =         127'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000; // D (0x00000010000000000000000000000020) 
14'h110e : LOC =         127'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000; // D (0x00000020000000000000000000000020) 
14'h17d2 : LOC =         127'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000; // D (0x00000040000000000000000000000020) 
14'h1a6a : LOC =         127'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000; // D (0x00000080000000000000000000000020) 
14'h011a : LOC =         127'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000; // D (0x00000100000000000000000000000020) 
14'h37fa : LOC =         127'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000; // D (0x00000200000000000000000000000020) 
14'h194d : LOC =         127'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000; // D (0x00000400000000000000000000000020) 
14'h0754 : LOC =         127'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000; // D (0x00000800000000000000000000000020) 
14'h3b66 : LOC =         127'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000; // D (0x00001000000000000000000000000020) 
14'h0075 : LOC =         127'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000; // D (0x00002000000000000000000000000020) 
14'h3524 : LOC =         127'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000; // D (0x00004000000000000000000000000020) 
14'h1cf1 : LOC =         127'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000; // D (0x00008000000000000000000000000020) 
14'h0c2c : LOC =         127'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000; // D (0x00010000000000000000000000000020) 
14'h2d96 : LOC =         127'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000; // D (0x00020000000000000000000000000020) 
14'h2d95 : LOC =         127'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000; // D (0x00040000000000000000000000000020) 
14'h2d93 : LOC =         127'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000; // D (0x00080000000000000000000000000020) 
14'h2d9f : LOC =         127'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000; // D (0x00100000000000000000000000000020) 
14'h2d87 : LOC =         127'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000; // D (0x00200000000000000000000000000020) 
14'h2db7 : LOC =         127'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000; // D (0x00400000000000000000000000000020) 
14'h2dd7 : LOC =         127'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000; // D (0x00800000000000000000000000000020) 
14'h2d17 : LOC =         127'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000; // D (0x01000000000000000000000000000020) 
14'h2c97 : LOC =         127'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000; // D (0x02000000000000000000000000000020) 
14'h2f97 : LOC =         127'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000; // D (0x04000000000000000000000000000020) 
14'h2997 : LOC =         127'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000; // D (0x08000000000000000000000000000020) 
14'h2597 : LOC =         127'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000; // D (0x10000000000000000000000000000020) 
14'h3d97 : LOC =         127'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000; // D (0x20000000000000000000000000000020) 
14'h0d97 : LOC =         127'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000; // D (0x40000000000000000000000000000020) 
14'h1859 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000; // S (0x00000000000000000000000000000040) 
14'h28eb : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000; // D (0x000000000000000000000000000000c0) 
14'h3a4a : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000000; // D (0x00000000000000000000000000000140) 
14'h1f08 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000; // D (0x00000000000000000000000000000240) 
14'h16fb : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000000; // D (0x00000000000000000000000000000440) 
14'h051d : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100001000000; // D (0x00000000000000000000000000000840) 
14'h22d1 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000001000000; // D (0x00000000000000000000000000001040) 
14'h2e3e : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000001000000; // D (0x00000000000000000000000000002040) 
14'h37e0 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000001000000; // D (0x00000000000000000000000000004040) 
14'h045c : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000001000000; // D (0x00000000000000000000000000008040) 
14'h2053 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000001000000; // D (0x00000000000000000000000000010040) 
14'h2b3a : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000001000000; // D (0x00000000000000000000000000020040) 
14'h3de8 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000001000000; // D (0x00000000000000000000000000040040) 
14'h104c : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000001000000; // D (0x00000000000000000000000000080040) 
14'h0873 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000001000000; // D (0x00000000000000000000000000100040) 
14'h380d : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000001000000; // D (0x00000000000000000000000000200040) 
14'h1b86 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001000000; // D (0x00000000000000000000000000400040) 
14'h1fe7 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000001000000; // D (0x00000000000000000000000000800040) 
14'h1725 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000001000000; // D (0x00000000000000000000000001000040) 
14'h06a1 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000001000000; // D (0x00000000000000000000000002000040) 
14'h25a9 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000001000000; // D (0x00000000000000000000000004000040) 
14'h20ce : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000001000000; // D (0x00000000000000000000000008000040) 
14'h2a00 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000001000000; // D (0x00000000000000000000000010000040) 
14'h3f9c : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000001000000; // D (0x00000000000000000000000020000040) 
14'h14a4 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000001000000; // D (0x00000000000000000000000040000040) 
14'h01a3 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000001000000; // D (0x00000000000000000000000080000040) 
14'h2bad : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000001000000; // D (0x00000000000000000000000100000040) 
14'h3cc6 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000001000000; // D (0x00000000000000000000000200000040) 
14'h1210 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000001000000; // D (0x00000000000000000000000400000040) 
14'h0ccb : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000001000000; // D (0x00000000000000000000000800000040) 
14'h317d : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000001000000; // D (0x00000000000000000000001000000040) 
14'h0966 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000001000000; // D (0x00000000000000000000002000000040) 
14'h3a27 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000001000000; // D (0x00000000000000000000004000000040) 
14'h1fd2 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000001000000; // D (0x00000000000000000000008000000040) 
14'h174f : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000001000000; // D (0x00000000000000000000010000000040) 
14'h0675 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000001000000; // D (0x00000000000000000000020000000040) 
14'h2401 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000001000000; // D (0x00000000000000000000040000000040) 
14'h239e : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000001000000; // D (0x00000000000000000000080000000040) 
14'h2ca0 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000; // D (0x00000000000000000000100000000040) 
14'h32dc : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000001000000; // D (0x00000000000000000000200000000040) 
14'h0e24 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000001000000; // D (0x00000000000000000000400000000040) 
14'h34a3 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000001000000; // D (0x00000000000000000000800000000040) 
14'h02da : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000001000000; // D (0x00000000000000000001000000000040) 
14'h2d5f : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000001000000; // D (0x00000000000000000002000000000040) 
14'h3122 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000001000000; // D (0x00000000000000000004000000000040) 
14'h09d8 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000001000000; // D (0x00000000000000000008000000000040) 
14'h3b5b : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000001000000; // D (0x00000000000000000010000000000040) 
14'h1d2a : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000001000000; // D (0x00000000000000000020000000000040) 
14'h12bf : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000001000000; // D (0x00000000000000000040000000000040) 
14'h0d95 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000001000000; // D (0x00000000000000000080000000000040) 
14'h33c1 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000001000000; // D (0x00000000000000000100000000000040) 
14'h0c1e : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000001000000; // D (0x00000000000000000200000000000040) 
14'h30d7 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000001000000; // D (0x00000000000000000400000000000040) 
14'h0a32 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000001000000; // D (0x00000000000000000800000000000040) 
14'h3c8f : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000001000000; // D (0x00000000000000001000000000000040) 
14'h1282 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000001000000; // D (0x00000000000000002000000000000040) 
14'h0def : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000001000000; // D (0x00000000000000004000000000000040) 
14'h3335 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000001000000; // D (0x00000000000000008000000000000040) 
14'h0df6 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000001000000; // D (0x00000000000000010000000000000040) 
14'h3307 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000001000000; // D (0x00000000000000020000000000000040) 
14'h0d92 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000001000000; // D (0x00000000000000040000000000000040) 
14'h33cf : LOC =         127'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000001000000; // D (0x00000000000000080000000000000040) 
14'h0c02 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000001000000; // D (0x00000000000000100000000000000040) 
14'h30ef : LOC =         127'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000001000000; // D (0x00000000000000200000000000000040) 
14'h0a42 : LOC =         127'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000001000000; // D (0x00000000000000400000000000000040) 
14'h3c6f : LOC =         127'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000001000000; // D (0x00000000000000800000000000000040) 
14'h1342 : LOC =         127'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000001000000; // D (0x00000000000001000000000000000040) 
14'h0e6f : LOC =         127'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000001000000; // D (0x00000000000002000000000000000040) 
14'h3435 : LOC =         127'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000001000000; // D (0x00000000000004000000000000000040) 
14'h03f6 : LOC =         127'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000001000000; // D (0x00000000000008000000000000000040) 
14'h2f07 : LOC =         127'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000001000000; // D (0x00000000000010000000000000000040) 
14'h3592 : LOC =         127'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000001000000; // D (0x00000000000020000000000000000040) 
14'h00b8 : LOC =         127'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000001000000; // D (0x00000000000040000000000000000040) 
14'h299b : LOC =         127'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000001000000; // D (0x00000000000080000000000000000040) 
14'h38aa : LOC =         127'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000001000000; // D (0x00000000000100000000000000000040) 
14'h1ac8 : LOC =         127'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000001000000; // D (0x00000000000200000000000000000040) 
14'h1d7b : LOC =         127'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000001000000; // D (0x00000000000400000000000000000040) 
14'h121d : LOC =         127'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000001000000; // D (0x00000000000800000000000000000040) 
14'h0cd1 : LOC =         127'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000001000000; // D (0x00000000001000000000000000000040) 
14'h3149 : LOC =         127'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000001000000; // D (0x00000000002000000000000000000040) 
14'h090e : LOC =         127'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000001000000; // D (0x00000000004000000000000000000040) 
14'h3af7 : LOC =         127'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000001000000; // D (0x00000000008000000000000000000040) 
14'h1e72 : LOC =         127'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000001000000; // D (0x00000000010000000000000000000040) 
14'h140f : LOC =         127'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000001000000; // D (0x00000000020000000000000000000040) 
14'h00f5 : LOC =         127'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000; // D (0x00000000040000000000000000000040) 
14'h2901 : LOC =         127'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000; // D (0x00000000080000000000000000000040) 
14'h399e : LOC =         127'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000; // D (0x00000000100000000000000000000040) 
14'h18a0 : LOC =         127'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000; // D (0x00000000200000000000000000000040) 
14'h19ab : LOC =         127'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000; // D (0x00000000400000000000000000000040) 
14'h1bbd : LOC =         127'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000; // D (0x00000000800000000000000000000040) 
14'h1f91 : LOC =         127'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000; // D (0x00000001000000000000000000000040) 
14'h17c9 : LOC =         127'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000; // D (0x00000002000000000000000000000040) 
14'h0779 : LOC =         127'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000; // D (0x00000004000000000000000000000040) 
14'h2619 : LOC =         127'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000; // D (0x00000008000000000000000000000040) 
14'h27ae : LOC =         127'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000; // D (0x00000010000000000000000000000040) 
14'h24c0 : LOC =         127'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000; // D (0x00000020000000000000000000000040) 
14'h221c : LOC =         127'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000; // D (0x00000040000000000000000000000040) 
14'h2fa4 : LOC =         127'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000; // D (0x00000080000000000000000000000040) 
14'h34d4 : LOC =         127'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000; // D (0x00000100000000000000000000000040) 
14'h0234 : LOC =         127'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000; // D (0x00000200000000000000000000000040) 
14'h2c83 : LOC =         127'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000; // D (0x00000400000000000000000000000040) 
14'h329a : LOC =         127'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000; // D (0x00000800000000000000000000000040) 
14'h0ea8 : LOC =         127'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000; // D (0x00001000000000000000000000000040) 
14'h35bb : LOC =         127'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000; // D (0x00002000000000000000000000000040) 
14'h00ea : LOC =         127'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000; // D (0x00004000000000000000000000000040) 
14'h293f : LOC =         127'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000; // D (0x00008000000000000000000000000040) 
14'h39e2 : LOC =         127'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000; // D (0x00010000000000000000000000000040) 
14'h1858 : LOC =         127'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000; // D (0x00020000000000000000000000000040) 
14'h185b : LOC =         127'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000; // D (0x00040000000000000000000000000040) 
14'h185d : LOC =         127'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000; // D (0x00080000000000000000000000000040) 
14'h1851 : LOC =         127'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000; // D (0x00100000000000000000000000000040) 
14'h1849 : LOC =         127'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000; // D (0x00200000000000000000000000000040) 
14'h1879 : LOC =         127'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000; // D (0x00400000000000000000000000000040) 
14'h1819 : LOC =         127'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000; // D (0x00800000000000000000000000000040) 
14'h18d9 : LOC =         127'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000; // D (0x01000000000000000000000000000040) 
14'h1959 : LOC =         127'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000; // D (0x02000000000000000000000000000040) 
14'h1a59 : LOC =         127'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000; // D (0x04000000000000000000000000000040) 
14'h1c59 : LOC =         127'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000; // D (0x08000000000000000000000000000040) 
14'h1059 : LOC =         127'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000; // D (0x10000000000000000000000000000040) 
14'h0859 : LOC =         127'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000; // D (0x20000000000000000000000000000040) 
14'h3859 : LOC =         127'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000; // D (0x40000000000000000000000000000040) 
14'h30b2 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000; // S (0x00000000000000000000000000000080) 
14'h12a1 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000; // D (0x00000000000000000000000000000180) 
14'h37e3 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000000; // D (0x00000000000000000000000000000280) 
14'h3e10 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000; // D (0x00000000000000000000000000000480) 
14'h2df6 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010000000; // D (0x00000000000000000000000000000880) 
14'h0a3a : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000010000000; // D (0x00000000000000000000000000001080) 
14'h06d5 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000010000000; // D (0x00000000000000000000000000002080) 
14'h1f0b : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000010000000; // D (0x00000000000000000000000000004080) 
14'h2cb7 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000010000000; // D (0x00000000000000000000000000008080) 
14'h08b8 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000010000000; // D (0x00000000000000000000000000010080) 
14'h03d1 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000010000000; // D (0x00000000000000000000000000020080) 
14'h1503 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000010000000; // D (0x00000000000000000000000000040080) 
14'h38a7 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000010000000; // D (0x00000000000000000000000000080080) 
14'h2098 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000010000000; // D (0x00000000000000000000000000100080) 
14'h10e6 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000010000000; // D (0x00000000000000000000000000200080) 
14'h336d : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000010000000; // D (0x00000000000000000000000000400080) 
14'h370c : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000010000000; // D (0x00000000000000000000000000800080) 
14'h3fce : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000010000000; // D (0x00000000000000000000000001000080) 
14'h2e4a : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000010000000; // D (0x00000000000000000000000002000080) 
14'h0d42 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000010000000; // D (0x00000000000000000000000004000080) 
14'h0825 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000010000000; // D (0x00000000000000000000000008000080) 
14'h02eb : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000010000000; // D (0x00000000000000000000000010000080) 
14'h1777 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000010000000; // D (0x00000000000000000000000020000080) 
14'h3c4f : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000010000000; // D (0x00000000000000000000000040000080) 
14'h2948 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000010000000; // D (0x00000000000000000000000080000080) 
14'h0346 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000010000000; // D (0x00000000000000000000000100000080) 
14'h142d : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000010000000; // D (0x00000000000000000000000200000080) 
14'h3afb : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000010000000; // D (0x00000000000000000000000400000080) 
14'h2420 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000010000000; // D (0x00000000000000000000000800000080) 
14'h1996 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000010000000; // D (0x00000000000000000000001000000080) 
14'h218d : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000010000000; // D (0x00000000000000000000002000000080) 
14'h12cc : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000010000000; // D (0x00000000000000000000004000000080) 
14'h3739 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000010000000; // D (0x00000000000000000000008000000080) 
14'h3fa4 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000010000000; // D (0x00000000000000000000010000000080) 
14'h2e9e : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000010000000; // D (0x00000000000000000000020000000080) 
14'h0cea : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000010000000; // D (0x00000000000000000000040000000080) 
14'h0b75 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000010000000; // D (0x00000000000000000000080000000080) 
14'h044b : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000010000000; // D (0x00000000000000000000100000000080) 
14'h1a37 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000010000000; // D (0x00000000000000000000200000000080) 
14'h26cf : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000010000000; // D (0x00000000000000000000400000000080) 
14'h1c48 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000010000000; // D (0x00000000000000000000800000000080) 
14'h2a31 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000010000000; // D (0x00000000000000000001000000000080) 
14'h05b4 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000010000000; // D (0x00000000000000000002000000000080) 
14'h19c9 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000010000000; // D (0x00000000000000000004000000000080) 
14'h2133 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000010000000; // D (0x00000000000000000008000000000080) 
14'h13b0 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000010000000; // D (0x00000000000000000010000000000080) 
14'h35c1 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000010000000; // D (0x00000000000000000020000000000080) 
14'h3a54 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000010000000; // D (0x00000000000000000040000000000080) 
14'h257e : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000010000000; // D (0x00000000000000000080000000000080) 
14'h1b2a : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000010000000; // D (0x00000000000000000100000000000080) 
14'h24f5 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000010000000; // D (0x00000000000000000200000000000080) 
14'h183c : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000010000000; // D (0x00000000000000000400000000000080) 
14'h22d9 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000010000000; // D (0x00000000000000000800000000000080) 
14'h1464 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000010000000; // D (0x00000000000000001000000000000080) 
14'h3a69 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000010000000; // D (0x00000000000000002000000000000080) 
14'h2504 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000010000000; // D (0x00000000000000004000000000000080) 
14'h1bde : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000010000000; // D (0x00000000000000008000000000000080) 
14'h251d : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000010000000; // D (0x00000000000000010000000000000080) 
14'h1bec : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000010000000; // D (0x00000000000000020000000000000080) 
14'h2579 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000010000000; // D (0x00000000000000040000000000000080) 
14'h1b24 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000010000000; // D (0x00000000000000080000000000000080) 
14'h24e9 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000010000000; // D (0x00000000000000100000000000000080) 
14'h1804 : LOC =         127'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000010000000; // D (0x00000000000000200000000000000080) 
14'h22a9 : LOC =         127'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000010000000; // D (0x00000000000000400000000000000080) 
14'h1484 : LOC =         127'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000010000000; // D (0x00000000000000800000000000000080) 
14'h3ba9 : LOC =         127'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000010000000; // D (0x00000000000001000000000000000080) 
14'h2684 : LOC =         127'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000010000000; // D (0x00000000000002000000000000000080) 
14'h1cde : LOC =         127'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000010000000; // D (0x00000000000004000000000000000080) 
14'h2b1d : LOC =         127'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000010000000; // D (0x00000000000008000000000000000080) 
14'h07ec : LOC =         127'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000010000000; // D (0x00000000000010000000000000000080) 
14'h1d79 : LOC =         127'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000010000000; // D (0x00000000000020000000000000000080) 
14'h2853 : LOC =         127'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000010000000; // D (0x00000000000040000000000000000080) 
14'h0170 : LOC =         127'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000010000000; // D (0x00000000000080000000000000000080) 
14'h1041 : LOC =         127'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000010000000; // D (0x00000000000100000000000000000080) 
14'h3223 : LOC =         127'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000010000000; // D (0x00000000000200000000000000000080) 
14'h3590 : LOC =         127'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000010000000; // D (0x00000000000400000000000000000080) 
14'h3af6 : LOC =         127'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000010000000; // D (0x00000000000800000000000000000080) 
14'h243a : LOC =         127'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000010000000; // D (0x00000000001000000000000000000080) 
14'h19a2 : LOC =         127'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000010000000; // D (0x00000000002000000000000000000080) 
14'h21e5 : LOC =         127'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000010000000; // D (0x00000000004000000000000000000080) 
14'h121c : LOC =         127'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000010000000; // D (0x00000000008000000000000000000080) 
14'h3699 : LOC =         127'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000010000000; // D (0x00000000010000000000000000000080) 
14'h3ce4 : LOC =         127'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000010000000; // D (0x00000000020000000000000000000080) 
14'h281e : LOC =         127'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000; // D (0x00000000040000000000000000000080) 
14'h01ea : LOC =         127'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000; // D (0x00000000080000000000000000000080) 
14'h1175 : LOC =         127'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000; // D (0x00000000100000000000000000000080) 
14'h304b : LOC =         127'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000; // D (0x00000000200000000000000000000080) 
14'h3140 : LOC =         127'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000; // D (0x00000000400000000000000000000080) 
14'h3356 : LOC =         127'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000; // D (0x00000000800000000000000000000080) 
14'h377a : LOC =         127'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000; // D (0x00000001000000000000000000000080) 
14'h3f22 : LOC =         127'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000; // D (0x00000002000000000000000000000080) 
14'h2f92 : LOC =         127'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000; // D (0x00000004000000000000000000000080) 
14'h0ef2 : LOC =         127'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000; // D (0x00000008000000000000000000000080) 
14'h0f45 : LOC =         127'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000; // D (0x00000010000000000000000000000080) 
14'h0c2b : LOC =         127'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000; // D (0x00000020000000000000000000000080) 
14'h0af7 : LOC =         127'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000; // D (0x00000040000000000000000000000080) 
14'h074f : LOC =         127'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000; // D (0x00000080000000000000000000000080) 
14'h1c3f : LOC =         127'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000; // D (0x00000100000000000000000000000080) 
14'h2adf : LOC =         127'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000; // D (0x00000200000000000000000000000080) 
14'h0468 : LOC =         127'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000; // D (0x00000400000000000000000000000080) 
14'h1a71 : LOC =         127'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000; // D (0x00000800000000000000000000000080) 
14'h2643 : LOC =         127'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000; // D (0x00001000000000000000000000000080) 
14'h1d50 : LOC =         127'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000; // D (0x00002000000000000000000000000080) 
14'h2801 : LOC =         127'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000; // D (0x00004000000000000000000000000080) 
14'h01d4 : LOC =         127'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000; // D (0x00008000000000000000000000000080) 
14'h1109 : LOC =         127'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000; // D (0x00010000000000000000000000000080) 
14'h30b3 : LOC =         127'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000; // D (0x00020000000000000000000000000080) 
14'h30b0 : LOC =         127'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000; // D (0x00040000000000000000000000000080) 
14'h30b6 : LOC =         127'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000; // D (0x00080000000000000000000000000080) 
14'h30ba : LOC =         127'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000; // D (0x00100000000000000000000000000080) 
14'h30a2 : LOC =         127'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000; // D (0x00200000000000000000000000000080) 
14'h3092 : LOC =         127'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000; // D (0x00400000000000000000000000000080) 
14'h30f2 : LOC =         127'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000; // D (0x00800000000000000000000000000080) 
14'h3032 : LOC =         127'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000; // D (0x01000000000000000000000000000080) 
14'h31b2 : LOC =         127'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000; // D (0x02000000000000000000000000000080) 
14'h32b2 : LOC =         127'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000; // D (0x04000000000000000000000000000080) 
14'h34b2 : LOC =         127'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000; // D (0x08000000000000000000000000000080) 
14'h38b2 : LOC =         127'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000; // D (0x10000000000000000000000000000080) 
14'h20b2 : LOC =         127'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000; // D (0x20000000000000000000000000000080) 
14'h10b2 : LOC =         127'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000; // D (0x40000000000000000000000000000080) 
14'h2213 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000; // S (0x00000000000000000000000000000100) 
14'h2542 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000; // D (0x00000000000000000000000000000300) 
14'h2cb1 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000; // D (0x00000000000000000000000000000500) 
14'h3f57 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000; // D (0x00000000000000000000000000000900) 
14'h189b : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000100000000; // D (0x00000000000000000000000000001100) 
14'h1474 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000100000000; // D (0x00000000000000000000000000002100) 
14'h0daa : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000100000000; // D (0x00000000000000000000000000004100) 
14'h3e16 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000100000000; // D (0x00000000000000000000000000008100) 
14'h1a19 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000100000000; // D (0x00000000000000000000000000010100) 
14'h1170 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000100000000; // D (0x00000000000000000000000000020100) 
14'h07a2 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000100000000; // D (0x00000000000000000000000000040100) 
14'h2a06 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000100000000; // D (0x00000000000000000000000000080100) 
14'h3239 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000100000000; // D (0x00000000000000000000000000100100) 
14'h0247 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000100000000; // D (0x00000000000000000000000000200100) 
14'h21cc : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000100000000; // D (0x00000000000000000000000000400100) 
14'h25ad : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000100000000; // D (0x00000000000000000000000000800100) 
14'h2d6f : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000100000000; // D (0x00000000000000000000000001000100) 
14'h3ceb : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000100000000; // D (0x00000000000000000000000002000100) 
14'h1fe3 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000100000000; // D (0x00000000000000000000000004000100) 
14'h1a84 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000100000000; // D (0x00000000000000000000000008000100) 
14'h104a : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000100000000; // D (0x00000000000000000000000010000100) 
14'h05d6 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000100000000; // D (0x00000000000000000000000020000100) 
14'h2eee : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000100000000; // D (0x00000000000000000000000040000100) 
14'h3be9 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000100000000; // D (0x00000000000000000000000080000100) 
14'h11e7 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000100000000; // D (0x00000000000000000000000100000100) 
14'h068c : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000100000000; // D (0x00000000000000000000000200000100) 
14'h285a : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000100000000; // D (0x00000000000000000000000400000100) 
14'h3681 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000100000000; // D (0x00000000000000000000000800000100) 
14'h0b37 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000100000000; // D (0x00000000000000000000001000000100) 
14'h332c : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000100000000; // D (0x00000000000000000000002000000100) 
14'h006d : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000100000000; // D (0x00000000000000000000004000000100) 
14'h2598 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000100000000; // D (0x00000000000000000000008000000100) 
14'h2d05 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000100000000; // D (0x00000000000000000000010000000100) 
14'h3c3f : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000100000000; // D (0x00000000000000000000020000000100) 
14'h1e4b : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000100000000; // D (0x00000000000000000000040000000100) 
14'h19d4 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000100000000; // D (0x00000000000000000000080000000100) 
14'h16ea : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000100000000; // D (0x00000000000000000000100000000100) 
14'h0896 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000100000000; // D (0x00000000000000000000200000000100) 
14'h346e : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000100000000; // D (0x00000000000000000000400000000100) 
14'h0ee9 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000100000000; // D (0x00000000000000000000800000000100) 
14'h3890 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000100000000; // D (0x00000000000000000001000000000100) 
14'h1715 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000100000000; // D (0x00000000000000000002000000000100) 
14'h0b68 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000100000000; // D (0x00000000000000000004000000000100) 
14'h3392 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000100000000; // D (0x00000000000000000008000000000100) 
14'h0111 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000100000000; // D (0x00000000000000000010000000000100) 
14'h2760 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000100000000; // D (0x00000000000000000020000000000100) 
14'h28f5 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000100000000; // D (0x00000000000000000040000000000100) 
14'h37df : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000100000000; // D (0x00000000000000000080000000000100) 
14'h098b : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000100000000; // D (0x00000000000000000100000000000100) 
14'h3654 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000100000000; // D (0x00000000000000000200000000000100) 
14'h0a9d : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000100000000; // D (0x00000000000000000400000000000100) 
14'h3078 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000100000000; // D (0x00000000000000000800000000000100) 
14'h06c5 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000100000000; // D (0x00000000000000001000000000000100) 
14'h28c8 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000100000000; // D (0x00000000000000002000000000000100) 
14'h37a5 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000100000000; // D (0x00000000000000004000000000000100) 
14'h097f : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000100000000; // D (0x00000000000000008000000000000100) 
14'h37bc : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000100000000; // D (0x00000000000000010000000000000100) 
14'h094d : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000100000000; // D (0x00000000000000020000000000000100) 
14'h37d8 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000100000000; // D (0x00000000000000040000000000000100) 
14'h0985 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000100000000; // D (0x00000000000000080000000000000100) 
14'h3648 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000100000000; // D (0x00000000000000100000000000000100) 
14'h0aa5 : LOC =         127'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000100000000; // D (0x00000000000000200000000000000100) 
14'h3008 : LOC =         127'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000100000000; // D (0x00000000000000400000000000000100) 
14'h0625 : LOC =         127'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000100000000; // D (0x00000000000000800000000000000100) 
14'h2908 : LOC =         127'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000100000000; // D (0x00000000000001000000000000000100) 
14'h3425 : LOC =         127'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000100000000; // D (0x00000000000002000000000000000100) 
14'h0e7f : LOC =         127'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000100000000; // D (0x00000000000004000000000000000100) 
14'h39bc : LOC =         127'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000100000000; // D (0x00000000000008000000000000000100) 
14'h154d : LOC =         127'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000100000000; // D (0x00000000000010000000000000000100) 
14'h0fd8 : LOC =         127'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000100000000; // D (0x00000000000020000000000000000100) 
14'h3af2 : LOC =         127'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000100000000; // D (0x00000000000040000000000000000100) 
14'h13d1 : LOC =         127'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000100000000; // D (0x00000000000080000000000000000100) 
14'h02e0 : LOC =         127'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000100000000; // D (0x00000000000100000000000000000100) 
14'h2082 : LOC =         127'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000100000000; // D (0x00000000000200000000000000000100) 
14'h2731 : LOC =         127'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000100000000; // D (0x00000000000400000000000000000100) 
14'h2857 : LOC =         127'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000100000000; // D (0x00000000000800000000000000000100) 
14'h369b : LOC =         127'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000100000000; // D (0x00000000001000000000000000000100) 
14'h0b03 : LOC =         127'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000100000000; // D (0x00000000002000000000000000000100) 
14'h3344 : LOC =         127'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000100000000; // D (0x00000000004000000000000000000100) 
14'h00bd : LOC =         127'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000100000000; // D (0x00000000008000000000000000000100) 
14'h2438 : LOC =         127'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000100000000; // D (0x00000000010000000000000000000100) 
14'h2e45 : LOC =         127'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000100000000; // D (0x00000000020000000000000000000100) 
14'h3abf : LOC =         127'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000; // D (0x00000000040000000000000000000100) 
14'h134b : LOC =         127'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000; // D (0x00000000080000000000000000000100) 
14'h03d4 : LOC =         127'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000; // D (0x00000000100000000000000000000100) 
14'h22ea : LOC =         127'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000; // D (0x00000000200000000000000000000100) 
14'h23e1 : LOC =         127'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000; // D (0x00000000400000000000000000000100) 
14'h21f7 : LOC =         127'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000; // D (0x00000000800000000000000000000100) 
14'h25db : LOC =         127'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000; // D (0x00000001000000000000000000000100) 
14'h2d83 : LOC =         127'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000; // D (0x00000002000000000000000000000100) 
14'h3d33 : LOC =         127'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000; // D (0x00000004000000000000000000000100) 
14'h1c53 : LOC =         127'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000; // D (0x00000008000000000000000000000100) 
14'h1de4 : LOC =         127'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000; // D (0x00000010000000000000000000000100) 
14'h1e8a : LOC =         127'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000; // D (0x00000020000000000000000000000100) 
14'h1856 : LOC =         127'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000; // D (0x00000040000000000000000000000100) 
14'h15ee : LOC =         127'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000; // D (0x00000080000000000000000000000100) 
14'h0e9e : LOC =         127'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000; // D (0x00000100000000000000000000000100) 
14'h387e : LOC =         127'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000; // D (0x00000200000000000000000000000100) 
14'h16c9 : LOC =         127'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000; // D (0x00000400000000000000000000000100) 
14'h08d0 : LOC =         127'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000; // D (0x00000800000000000000000000000100) 
14'h34e2 : LOC =         127'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000; // D (0x00001000000000000000000000000100) 
14'h0ff1 : LOC =         127'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000; // D (0x00002000000000000000000000000100) 
14'h3aa0 : LOC =         127'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000; // D (0x00004000000000000000000000000100) 
14'h1375 : LOC =         127'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000; // D (0x00008000000000000000000000000100) 
14'h03a8 : LOC =         127'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000; // D (0x00010000000000000000000000000100) 
14'h2212 : LOC =         127'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000; // D (0x00020000000000000000000000000100) 
14'h2211 : LOC =         127'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000; // D (0x00040000000000000000000000000100) 
14'h2217 : LOC =         127'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000; // D (0x00080000000000000000000000000100) 
14'h221b : LOC =         127'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000; // D (0x00100000000000000000000000000100) 
14'h2203 : LOC =         127'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000; // D (0x00200000000000000000000000000100) 
14'h2233 : LOC =         127'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000; // D (0x00400000000000000000000000000100) 
14'h2253 : LOC =         127'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000; // D (0x00800000000000000000000000000100) 
14'h2293 : LOC =         127'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000; // D (0x01000000000000000000000000000100) 
14'h2313 : LOC =         127'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000; // D (0x02000000000000000000000000000100) 
14'h2013 : LOC =         127'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000; // D (0x04000000000000000000000000000100) 
14'h2613 : LOC =         127'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000; // D (0x08000000000000000000000000000100) 
14'h2a13 : LOC =         127'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000; // D (0x10000000000000000000000000000100) 
14'h3213 : LOC =         127'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000; // D (0x20000000000000000000000000000100) 
14'h0213 : LOC =         127'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000; // D (0x40000000000000000000000000000100) 
14'h0751 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000; // S (0x00000000000000000000000000000200) 
14'h09f3 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000; // D (0x00000000000000000000000000000600) 
14'h1a15 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000000000; // D (0x00000000000000000000000000000a00) 
14'h3dd9 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000000; // D (0x00000000000000000000000000001200) 
14'h3136 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000000000; // D (0x00000000000000000000000000002200) 
14'h28e8 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100001000000000; // D (0x00000000000000000000000000004200) 
14'h1b54 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000001000000000; // D (0x00000000000000000000000000008200) 
14'h3f5b : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000001000000000; // D (0x00000000000000000000000000010200) 
14'h3432 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000001000000000; // D (0x00000000000000000000000000020200) 
14'h22e0 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000001000000000; // D (0x00000000000000000000000000040200) 
14'h0f44 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000001000000000; // D (0x00000000000000000000000000080200) 
14'h177b : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000001000000000; // D (0x00000000000000000000000000100200) 
14'h2705 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000001000000000; // D (0x00000000000000000000000000200200) 
14'h048e : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000001000000000; // D (0x00000000000000000000000000400200) 
14'h00ef : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000001000000000; // D (0x00000000000000000000000000800200) 
14'h082d : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000001000000000; // D (0x00000000000000000000000001000200) 
14'h19a9 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001000000000; // D (0x00000000000000000000000002000200) 
14'h3aa1 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000001000000000; // D (0x00000000000000000000000004000200) 
14'h3fc6 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000001000000000; // D (0x00000000000000000000000008000200) 
14'h3508 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000001000000000; // D (0x00000000000000000000000010000200) 
14'h2094 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000001000000000; // D (0x00000000000000000000000020000200) 
14'h0bac : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000001000000000; // D (0x00000000000000000000000040000200) 
14'h1eab : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000001000000000; // D (0x00000000000000000000000080000200) 
14'h34a5 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000001000000000; // D (0x00000000000000000000000100000200) 
14'h23ce : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000001000000000; // D (0x00000000000000000000000200000200) 
14'h0d18 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000001000000000; // D (0x00000000000000000000000400000200) 
14'h13c3 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000001000000000; // D (0x00000000000000000000000800000200) 
14'h2e75 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000001000000000; // D (0x00000000000000000000001000000200) 
14'h166e : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000001000000000; // D (0x00000000000000000000002000000200) 
14'h252f : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000001000000000; // D (0x00000000000000000000004000000200) 
14'h00da : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000001000000000; // D (0x00000000000000000000008000000200) 
14'h0847 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000001000000000; // D (0x00000000000000000000010000000200) 
14'h197d : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000001000000000; // D (0x00000000000000000000020000000200) 
14'h3b09 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000001000000000; // D (0x00000000000000000000040000000200) 
14'h3c96 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000001000000000; // D (0x00000000000000000000080000000200) 
14'h33a8 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000001000000000; // D (0x00000000000000000000100000000200) 
14'h2dd4 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000001000000000; // D (0x00000000000000000000200000000200) 
14'h112c : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000001000000000; // D (0x00000000000000000000400000000200) 
14'h2bab : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000; // D (0x00000000000000000000800000000200) 
14'h1dd2 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000001000000000; // D (0x00000000000000000001000000000200) 
14'h3257 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000001000000000; // D (0x00000000000000000002000000000200) 
14'h2e2a : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000001000000000; // D (0x00000000000000000004000000000200) 
14'h16d0 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000001000000000; // D (0x00000000000000000008000000000200) 
14'h2453 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000001000000000; // D (0x00000000000000000010000000000200) 
14'h0222 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000001000000000; // D (0x00000000000000000020000000000200) 
14'h0db7 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000001000000000; // D (0x00000000000000000040000000000200) 
14'h129d : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000001000000000; // D (0x00000000000000000080000000000200) 
14'h2cc9 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000001000000000; // D (0x00000000000000000100000000000200) 
14'h1316 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000001000000000; // D (0x00000000000000000200000000000200) 
14'h2fdf : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000001000000000; // D (0x00000000000000000400000000000200) 
14'h153a : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000001000000000; // D (0x00000000000000000800000000000200) 
14'h2387 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000001000000000; // D (0x00000000000000001000000000000200) 
14'h0d8a : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000001000000000; // D (0x00000000000000002000000000000200) 
14'h12e7 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000001000000000; // D (0x00000000000000004000000000000200) 
14'h2c3d : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000001000000000; // D (0x00000000000000008000000000000200) 
14'h12fe : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000001000000000; // D (0x00000000000000010000000000000200) 
14'h2c0f : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000001000000000; // D (0x00000000000000020000000000000200) 
14'h129a : LOC =         127'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000001000000000; // D (0x00000000000000040000000000000200) 
14'h2cc7 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000001000000000; // D (0x00000000000000080000000000000200) 
14'h130a : LOC =         127'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000001000000000; // D (0x00000000000000100000000000000200) 
14'h2fe7 : LOC =         127'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000001000000000; // D (0x00000000000000200000000000000200) 
14'h154a : LOC =         127'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000001000000000; // D (0x00000000000000400000000000000200) 
14'h2367 : LOC =         127'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000001000000000; // D (0x00000000000000800000000000000200) 
14'h0c4a : LOC =         127'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000001000000000; // D (0x00000000000001000000000000000200) 
14'h1167 : LOC =         127'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000001000000000; // D (0x00000000000002000000000000000200) 
14'h2b3d : LOC =         127'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000001000000000; // D (0x00000000000004000000000000000200) 
14'h1cfe : LOC =         127'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000001000000000; // D (0x00000000000008000000000000000200) 
14'h300f : LOC =         127'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000001000000000; // D (0x00000000000010000000000000000200) 
14'h2a9a : LOC =         127'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000001000000000; // D (0x00000000000020000000000000000200) 
14'h1fb0 : LOC =         127'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000001000000000; // D (0x00000000000040000000000000000200) 
14'h3693 : LOC =         127'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000001000000000; // D (0x00000000000080000000000000000200) 
14'h27a2 : LOC =         127'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000001000000000; // D (0x00000000000100000000000000000200) 
14'h05c0 : LOC =         127'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000001000000000; // D (0x00000000000200000000000000000200) 
14'h0273 : LOC =         127'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000001000000000; // D (0x00000000000400000000000000000200) 
14'h0d15 : LOC =         127'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000001000000000; // D (0x00000000000800000000000000000200) 
14'h13d9 : LOC =         127'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000001000000000; // D (0x00000000001000000000000000000200) 
14'h2e41 : LOC =         127'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000001000000000; // D (0x00000000002000000000000000000200) 
14'h1606 : LOC =         127'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000001000000000; // D (0x00000000004000000000000000000200) 
14'h25ff : LOC =         127'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000001000000000; // D (0x00000000008000000000000000000200) 
14'h017a : LOC =         127'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000001000000000; // D (0x00000000010000000000000000000200) 
14'h0b07 : LOC =         127'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000001000000000; // D (0x00000000020000000000000000000200) 
14'h1ffd : LOC =         127'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000; // D (0x00000000040000000000000000000200) 
14'h3609 : LOC =         127'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000; // D (0x00000000080000000000000000000200) 
14'h2696 : LOC =         127'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000; // D (0x00000000100000000000000000000200) 
14'h07a8 : LOC =         127'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000; // D (0x00000000200000000000000000000200) 
14'h06a3 : LOC =         127'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000; // D (0x00000000400000000000000000000200) 
14'h04b5 : LOC =         127'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000; // D (0x00000000800000000000000000000200) 
14'h0099 : LOC =         127'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000; // D (0x00000001000000000000000000000200) 
14'h08c1 : LOC =         127'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000; // D (0x00000002000000000000000000000200) 
14'h1871 : LOC =         127'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000; // D (0x00000004000000000000000000000200) 
14'h3911 : LOC =         127'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000; // D (0x00000008000000000000000000000200) 
14'h38a6 : LOC =         127'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000; // D (0x00000010000000000000000000000200) 
14'h3bc8 : LOC =         127'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000; // D (0x00000020000000000000000000000200) 
14'h3d14 : LOC =         127'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000; // D (0x00000040000000000000000000000200) 
14'h30ac : LOC =         127'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000; // D (0x00000080000000000000000000000200) 
14'h2bdc : LOC =         127'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000; // D (0x00000100000000000000000000000200) 
14'h1d3c : LOC =         127'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000; // D (0x00000200000000000000000000000200) 
14'h338b : LOC =         127'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000; // D (0x00000400000000000000000000000200) 
14'h2d92 : LOC =         127'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000; // D (0x00000800000000000000000000000200) 
14'h11a0 : LOC =         127'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000; // D (0x00001000000000000000000000000200) 
14'h2ab3 : LOC =         127'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000; // D (0x00002000000000000000000000000200) 
14'h1fe2 : LOC =         127'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000; // D (0x00004000000000000000000000000200) 
14'h3637 : LOC =         127'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000; // D (0x00008000000000000000000000000200) 
14'h26ea : LOC =         127'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000; // D (0x00010000000000000000000000000200) 
14'h0750 : LOC =         127'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000; // D (0x00020000000000000000000000000200) 
14'h0753 : LOC =         127'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000; // D (0x00040000000000000000000000000200) 
14'h0755 : LOC =         127'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000; // D (0x00080000000000000000000000000200) 
14'h0759 : LOC =         127'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000; // D (0x00100000000000000000000000000200) 
14'h0741 : LOC =         127'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000; // D (0x00200000000000000000000000000200) 
14'h0771 : LOC =         127'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000; // D (0x00400000000000000000000000000200) 
14'h0711 : LOC =         127'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000; // D (0x00800000000000000000000000000200) 
14'h07d1 : LOC =         127'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000; // D (0x01000000000000000000000000000200) 
14'h0651 : LOC =         127'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000; // D (0x02000000000000000000000000000200) 
14'h0551 : LOC =         127'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000; // D (0x04000000000000000000000000000200) 
14'h0351 : LOC =         127'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000; // D (0x08000000000000000000000000000200) 
14'h0f51 : LOC =         127'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000; // D (0x10000000000000000000000000000200) 
14'h1751 : LOC =         127'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000; // D (0x20000000000000000000000000000200) 
14'h2751 : LOC =         127'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000; // D (0x40000000000000000000000000000200) 
14'h0ea2 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000; // S (0x00000000000000000000000000000400) 
14'h13e6 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000; // D (0x00000000000000000000000000000c00) 
14'h342a : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000000000; // D (0x00000000000000000000000000001400) 
14'h38c5 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000; // D (0x00000000000000000000000000002400) 
14'h211b : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010000000000; // D (0x00000000000000000000000000004400) 
14'h12a7 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000010000000000; // D (0x00000000000000000000000000008400) 
14'h36a8 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000010000000000; // D (0x00000000000000000000000000010400) 
14'h3dc1 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000010000000000; // D (0x00000000000000000000000000020400) 
14'h2b13 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000010000000000; // D (0x00000000000000000000000000040400) 
14'h06b7 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000010000000000; // D (0x00000000000000000000000000080400) 
14'h1e88 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000010000000000; // D (0x00000000000000000000000000100400) 
14'h2ef6 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000010000000000; // D (0x00000000000000000000000000200400) 
14'h0d7d : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000010000000000; // D (0x00000000000000000000000000400400) 
14'h091c : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000010000000000; // D (0x00000000000000000000000000800400) 
14'h01de : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000010000000000; // D (0x00000000000000000000000001000400) 
14'h105a : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000010000000000; // D (0x00000000000000000000000002000400) 
14'h3352 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000010000000000; // D (0x00000000000000000000000004000400) 
14'h3635 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000010000000000; // D (0x00000000000000000000000008000400) 
14'h3cfb : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000010000000000; // D (0x00000000000000000000000010000400) 
14'h2967 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000010000000000; // D (0x00000000000000000000000020000400) 
14'h025f : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000010000000000; // D (0x00000000000000000000000040000400) 
14'h1758 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000010000000000; // D (0x00000000000000000000000080000400) 
14'h3d56 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000010000000000; // D (0x00000000000000000000000100000400) 
14'h2a3d : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000010000000000; // D (0x00000000000000000000000200000400) 
14'h04eb : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000010000000000; // D (0x00000000000000000000000400000400) 
14'h1a30 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000010000000000; // D (0x00000000000000000000000800000400) 
14'h2786 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000010000000000; // D (0x00000000000000000000001000000400) 
14'h1f9d : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000010000000000; // D (0x00000000000000000000002000000400) 
14'h2cdc : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000010000000000; // D (0x00000000000000000000004000000400) 
14'h0929 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000010000000000; // D (0x00000000000000000000008000000400) 
14'h01b4 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000010000000000; // D (0x00000000000000000000010000000400) 
14'h108e : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000010000000000; // D (0x00000000000000000000020000000400) 
14'h32fa : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000010000000000; // D (0x00000000000000000000040000000400) 
14'h3565 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000010000000000; // D (0x00000000000000000000080000000400) 
14'h3a5b : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000010000000000; // D (0x00000000000000000000100000000400) 
14'h2427 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000010000000000; // D (0x00000000000000000000200000000400) 
14'h18df : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000010000000000; // D (0x00000000000000000000400000000400) 
14'h2258 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000010000000000; // D (0x00000000000000000000800000000400) 
14'h1421 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000010000000000; // D (0x00000000000000000001000000000400) 
14'h3ba4 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000010000000000; // D (0x00000000000000000002000000000400) 
14'h27d9 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000010000000000; // D (0x00000000000000000004000000000400) 
14'h1f23 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000010000000000; // D (0x00000000000000000008000000000400) 
14'h2da0 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000010000000000; // D (0x00000000000000000010000000000400) 
14'h0bd1 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000010000000000; // D (0x00000000000000000020000000000400) 
14'h0444 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000010000000000; // D (0x00000000000000000040000000000400) 
14'h1b6e : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000010000000000; // D (0x00000000000000000080000000000400) 
14'h253a : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000010000000000; // D (0x00000000000000000100000000000400) 
14'h1ae5 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000010000000000; // D (0x00000000000000000200000000000400) 
14'h262c : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000010000000000; // D (0x00000000000000000400000000000400) 
14'h1cc9 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000010000000000; // D (0x00000000000000000800000000000400) 
14'h2a74 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000010000000000; // D (0x00000000000000001000000000000400) 
14'h0479 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000010000000000; // D (0x00000000000000002000000000000400) 
14'h1b14 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000010000000000; // D (0x00000000000000004000000000000400) 
14'h25ce : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000010000000000; // D (0x00000000000000008000000000000400) 
14'h1b0d : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000010000000000; // D (0x00000000000000010000000000000400) 
14'h25fc : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000010000000000; // D (0x00000000000000020000000000000400) 
14'h1b69 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000010000000000; // D (0x00000000000000040000000000000400) 
14'h2534 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000010000000000; // D (0x00000000000000080000000000000400) 
14'h1af9 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000010000000000; // D (0x00000000000000100000000000000400) 
14'h2614 : LOC =         127'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000010000000000; // D (0x00000000000000200000000000000400) 
14'h1cb9 : LOC =         127'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000010000000000; // D (0x00000000000000400000000000000400) 
14'h2a94 : LOC =         127'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000010000000000; // D (0x00000000000000800000000000000400) 
14'h05b9 : LOC =         127'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000010000000000; // D (0x00000000000001000000000000000400) 
14'h1894 : LOC =         127'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000010000000000; // D (0x00000000000002000000000000000400) 
14'h22ce : LOC =         127'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000010000000000; // D (0x00000000000004000000000000000400) 
14'h150d : LOC =         127'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000010000000000; // D (0x00000000000008000000000000000400) 
14'h39fc : LOC =         127'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000010000000000; // D (0x00000000000010000000000000000400) 
14'h2369 : LOC =         127'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000010000000000; // D (0x00000000000020000000000000000400) 
14'h1643 : LOC =         127'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000010000000000; // D (0x00000000000040000000000000000400) 
14'h3f60 : LOC =         127'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000010000000000; // D (0x00000000000080000000000000000400) 
14'h2e51 : LOC =         127'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000010000000000; // D (0x00000000000100000000000000000400) 
14'h0c33 : LOC =         127'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000010000000000; // D (0x00000000000200000000000000000400) 
14'h0b80 : LOC =         127'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000010000000000; // D (0x00000000000400000000000000000400) 
14'h04e6 : LOC =         127'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000010000000000; // D (0x00000000000800000000000000000400) 
14'h1a2a : LOC =         127'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000010000000000; // D (0x00000000001000000000000000000400) 
14'h27b2 : LOC =         127'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000010000000000; // D (0x00000000002000000000000000000400) 
14'h1ff5 : LOC =         127'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000010000000000; // D (0x00000000004000000000000000000400) 
14'h2c0c : LOC =         127'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000010000000000; // D (0x00000000008000000000000000000400) 
14'h0889 : LOC =         127'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000010000000000; // D (0x00000000010000000000000000000400) 
14'h02f4 : LOC =         127'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000010000000000; // D (0x00000000020000000000000000000400) 
14'h160e : LOC =         127'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000; // D (0x00000000040000000000000000000400) 
14'h3ffa : LOC =         127'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000; // D (0x00000000080000000000000000000400) 
14'h2f65 : LOC =         127'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000; // D (0x00000000100000000000000000000400) 
14'h0e5b : LOC =         127'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000; // D (0x00000000200000000000000000000400) 
14'h0f50 : LOC =         127'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000; // D (0x00000000400000000000000000000400) 
14'h0d46 : LOC =         127'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000; // D (0x00000000800000000000000000000400) 
14'h096a : LOC =         127'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000; // D (0x00000001000000000000000000000400) 
14'h0132 : LOC =         127'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000; // D (0x00000002000000000000000000000400) 
14'h1182 : LOC =         127'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000; // D (0x00000004000000000000000000000400) 
14'h30e2 : LOC =         127'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000; // D (0x00000008000000000000000000000400) 
14'h3155 : LOC =         127'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000; // D (0x00000010000000000000000000000400) 
14'h323b : LOC =         127'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000; // D (0x00000020000000000000000000000400) 
14'h34e7 : LOC =         127'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000; // D (0x00000040000000000000000000000400) 
14'h395f : LOC =         127'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000; // D (0x00000080000000000000000000000400) 
14'h222f : LOC =         127'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000; // D (0x00000100000000000000000000000400) 
14'h14cf : LOC =         127'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000; // D (0x00000200000000000000000000000400) 
14'h3a78 : LOC =         127'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000; // D (0x00000400000000000000000000000400) 
14'h2461 : LOC =         127'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000; // D (0x00000800000000000000000000000400) 
14'h1853 : LOC =         127'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000; // D (0x00001000000000000000000000000400) 
14'h2340 : LOC =         127'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000; // D (0x00002000000000000000000000000400) 
14'h1611 : LOC =         127'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000; // D (0x00004000000000000000000000000400) 
14'h3fc4 : LOC =         127'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000; // D (0x00008000000000000000000000000400) 
14'h2f19 : LOC =         127'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000; // D (0x00010000000000000000000000000400) 
14'h0ea3 : LOC =         127'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000; // D (0x00020000000000000000000000000400) 
14'h0ea0 : LOC =         127'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000; // D (0x00040000000000000000000000000400) 
14'h0ea6 : LOC =         127'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000; // D (0x00080000000000000000000000000400) 
14'h0eaa : LOC =         127'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000; // D (0x00100000000000000000000000000400) 
14'h0eb2 : LOC =         127'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000; // D (0x00200000000000000000000000000400) 
14'h0e82 : LOC =         127'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000; // D (0x00400000000000000000000000000400) 
14'h0ee2 : LOC =         127'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000; // D (0x00800000000000000000000000000400) 
14'h0e22 : LOC =         127'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000; // D (0x01000000000000000000000000000400) 
14'h0fa2 : LOC =         127'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000; // D (0x02000000000000000000000000000400) 
14'h0ca2 : LOC =         127'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000; // D (0x04000000000000000000000000000400) 
14'h0aa2 : LOC =         127'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000; // D (0x08000000000000000000000000000400) 
14'h06a2 : LOC =         127'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000; // D (0x10000000000000000000000000000400) 
14'h1ea2 : LOC =         127'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000; // D (0x20000000000000000000000000000400) 
14'h2ea2 : LOC =         127'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000; // D (0x40000000000000000000000000000400) 
14'h1d44 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000; // S (0x00000000000000000000000000000800) 
14'h27cc : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000; // D (0x00000000000000000000000000001800) 
14'h2b23 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000; // D (0x00000000000000000000000000002800) 
14'h32fd : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000; // D (0x00000000000000000000000000004800) 
14'h0141 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000100000000000; // D (0x00000000000000000000000000008800) 
14'h254e : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000100000000000; // D (0x00000000000000000000000000010800) 
14'h2e27 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000100000000000; // D (0x00000000000000000000000000020800) 
14'h38f5 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000100000000000; // D (0x00000000000000000000000000040800) 
14'h1551 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000100000000000; // D (0x00000000000000000000000000080800) 
14'h0d6e : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000100000000000; // D (0x00000000000000000000000000100800) 
14'h3d10 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000100000000000; // D (0x00000000000000000000000000200800) 
14'h1e9b : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000100000000000; // D (0x00000000000000000000000000400800) 
14'h1afa : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000100000000000; // D (0x00000000000000000000000000800800) 
14'h1238 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000100000000000; // D (0x00000000000000000000000001000800) 
14'h03bc : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000100000000000; // D (0x00000000000000000000000002000800) 
14'h20b4 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000100000000000; // D (0x00000000000000000000000004000800) 
14'h25d3 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000100000000000; // D (0x00000000000000000000000008000800) 
14'h2f1d : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000100000000000; // D (0x00000000000000000000000010000800) 
14'h3a81 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000100000000000; // D (0x00000000000000000000000020000800) 
14'h11b9 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000100000000000; // D (0x00000000000000000000000040000800) 
14'h04be : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000100000000000; // D (0x00000000000000000000000080000800) 
14'h2eb0 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000100000000000; // D (0x00000000000000000000000100000800) 
14'h39db : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000100000000000; // D (0x00000000000000000000000200000800) 
14'h170d : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000100000000000; // D (0x00000000000000000000000400000800) 
14'h09d6 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000100000000000; // D (0x00000000000000000000000800000800) 
14'h3460 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000100000000000; // D (0x00000000000000000000001000000800) 
14'h0c7b : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000100000000000; // D (0x00000000000000000000002000000800) 
14'h3f3a : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000100000000000; // D (0x00000000000000000000004000000800) 
14'h1acf : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000100000000000; // D (0x00000000000000000000008000000800) 
14'h1252 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000100000000000; // D (0x00000000000000000000010000000800) 
14'h0368 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000100000000000; // D (0x00000000000000000000020000000800) 
14'h211c : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000100000000000; // D (0x00000000000000000000040000000800) 
14'h2683 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000100000000000; // D (0x00000000000000000000080000000800) 
14'h29bd : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000100000000000; // D (0x00000000000000000000100000000800) 
14'h37c1 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000100000000000; // D (0x00000000000000000000200000000800) 
14'h0b39 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000100000000000; // D (0x00000000000000000000400000000800) 
14'h31be : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000100000000000; // D (0x00000000000000000000800000000800) 
14'h07c7 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000100000000000; // D (0x00000000000000000001000000000800) 
14'h2842 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000100000000000; // D (0x00000000000000000002000000000800) 
14'h343f : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000100000000000; // D (0x00000000000000000004000000000800) 
14'h0cc5 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000100000000000; // D (0x00000000000000000008000000000800) 
14'h3e46 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000100000000000; // D (0x00000000000000000010000000000800) 
14'h1837 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000100000000000; // D (0x00000000000000000020000000000800) 
14'h17a2 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000100000000000; // D (0x00000000000000000040000000000800) 
14'h0888 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000100000000000; // D (0x00000000000000000080000000000800) 
14'h36dc : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000100000000000; // D (0x00000000000000000100000000000800) 
14'h0903 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000100000000000; // D (0x00000000000000000200000000000800) 
14'h35ca : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000100000000000; // D (0x00000000000000000400000000000800) 
14'h0f2f : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000100000000000; // D (0x00000000000000000800000000000800) 
14'h3992 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000100000000000; // D (0x00000000000000001000000000000800) 
14'h179f : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000100000000000; // D (0x00000000000000002000000000000800) 
14'h08f2 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000100000000000; // D (0x00000000000000004000000000000800) 
14'h3628 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000100000000000; // D (0x00000000000000008000000000000800) 
14'h08eb : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000100000000000; // D (0x00000000000000010000000000000800) 
14'h361a : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000100000000000; // D (0x00000000000000020000000000000800) 
14'h088f : LOC =         127'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000100000000000; // D (0x00000000000000040000000000000800) 
14'h36d2 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000100000000000; // D (0x00000000000000080000000000000800) 
14'h091f : LOC =         127'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000100000000000; // D (0x00000000000000100000000000000800) 
14'h35f2 : LOC =         127'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000100000000000; // D (0x00000000000000200000000000000800) 
14'h0f5f : LOC =         127'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000100000000000; // D (0x00000000000000400000000000000800) 
14'h3972 : LOC =         127'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000100000000000; // D (0x00000000000000800000000000000800) 
14'h165f : LOC =         127'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000100000000000; // D (0x00000000000001000000000000000800) 
14'h0b72 : LOC =         127'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000100000000000; // D (0x00000000000002000000000000000800) 
14'h3128 : LOC =         127'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000100000000000; // D (0x00000000000004000000000000000800) 
14'h06eb : LOC =         127'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000100000000000; // D (0x00000000000008000000000000000800) 
14'h2a1a : LOC =         127'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000100000000000; // D (0x00000000000010000000000000000800) 
14'h308f : LOC =         127'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000100000000000; // D (0x00000000000020000000000000000800) 
14'h05a5 : LOC =         127'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000100000000000; // D (0x00000000000040000000000000000800) 
14'h2c86 : LOC =         127'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000100000000000; // D (0x00000000000080000000000000000800) 
14'h3db7 : LOC =         127'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000100000000000; // D (0x00000000000100000000000000000800) 
14'h1fd5 : LOC =         127'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000100000000000; // D (0x00000000000200000000000000000800) 
14'h1866 : LOC =         127'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000100000000000; // D (0x00000000000400000000000000000800) 
14'h1700 : LOC =         127'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000100000000000; // D (0x00000000000800000000000000000800) 
14'h09cc : LOC =         127'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000100000000000; // D (0x00000000001000000000000000000800) 
14'h3454 : LOC =         127'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000100000000000; // D (0x00000000002000000000000000000800) 
14'h0c13 : LOC =         127'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000100000000000; // D (0x00000000004000000000000000000800) 
14'h3fea : LOC =         127'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000100000000000; // D (0x00000000008000000000000000000800) 
14'h1b6f : LOC =         127'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000100000000000; // D (0x00000000010000000000000000000800) 
14'h1112 : LOC =         127'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000100000000000; // D (0x00000000020000000000000000000800) 
14'h05e8 : LOC =         127'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000; // D (0x00000000040000000000000000000800) 
14'h2c1c : LOC =         127'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000; // D (0x00000000080000000000000000000800) 
14'h3c83 : LOC =         127'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000; // D (0x00000000100000000000000000000800) 
14'h1dbd : LOC =         127'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000; // D (0x00000000200000000000000000000800) 
14'h1cb6 : LOC =         127'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000; // D (0x00000000400000000000000000000800) 
14'h1ea0 : LOC =         127'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000; // D (0x00000000800000000000000000000800) 
14'h1a8c : LOC =         127'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000; // D (0x00000001000000000000000000000800) 
14'h12d4 : LOC =         127'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000; // D (0x00000002000000000000000000000800) 
14'h0264 : LOC =         127'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000; // D (0x00000004000000000000000000000800) 
14'h2304 : LOC =         127'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000; // D (0x00000008000000000000000000000800) 
14'h22b3 : LOC =         127'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000; // D (0x00000010000000000000000000000800) 
14'h21dd : LOC =         127'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000; // D (0x00000020000000000000000000000800) 
14'h2701 : LOC =         127'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000; // D (0x00000040000000000000000000000800) 
14'h2ab9 : LOC =         127'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000; // D (0x00000080000000000000000000000800) 
14'h31c9 : LOC =         127'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000; // D (0x00000100000000000000000000000800) 
14'h0729 : LOC =         127'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000; // D (0x00000200000000000000000000000800) 
14'h299e : LOC =         127'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000; // D (0x00000400000000000000000000000800) 
14'h3787 : LOC =         127'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000; // D (0x00000800000000000000000000000800) 
14'h0bb5 : LOC =         127'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000; // D (0x00001000000000000000000000000800) 
14'h30a6 : LOC =         127'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000; // D (0x00002000000000000000000000000800) 
14'h05f7 : LOC =         127'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000; // D (0x00004000000000000000000000000800) 
14'h2c22 : LOC =         127'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000; // D (0x00008000000000000000000000000800) 
14'h3cff : LOC =         127'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000; // D (0x00010000000000000000000000000800) 
14'h1d45 : LOC =         127'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000; // D (0x00020000000000000000000000000800) 
14'h1d46 : LOC =         127'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000; // D (0x00040000000000000000000000000800) 
14'h1d40 : LOC =         127'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000; // D (0x00080000000000000000000000000800) 
14'h1d4c : LOC =         127'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000; // D (0x00100000000000000000000000000800) 
14'h1d54 : LOC =         127'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000; // D (0x00200000000000000000000000000800) 
14'h1d64 : LOC =         127'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000; // D (0x00400000000000000000000000000800) 
14'h1d04 : LOC =         127'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000; // D (0x00800000000000000000000000000800) 
14'h1dc4 : LOC =         127'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000; // D (0x01000000000000000000000000000800) 
14'h1c44 : LOC =         127'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000; // D (0x02000000000000000000000000000800) 
14'h1f44 : LOC =         127'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000; // D (0x04000000000000000000000000000800) 
14'h1944 : LOC =         127'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000; // D (0x08000000000000000000000000000800) 
14'h1544 : LOC =         127'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000; // D (0x10000000000000000000000000000800) 
14'h0d44 : LOC =         127'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000; // D (0x20000000000000000000000000000800) 
14'h3d44 : LOC =         127'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000; // D (0x40000000000000000000000000000800) 
14'h3a88 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000; // S (0x00000000000000000000000000001000) 
14'h0cef : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000; // D (0x00000000000000000000000000003000) 
14'h1531 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000000000000; // D (0x00000000000000000000000000005000) 
14'h268d : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000000000; // D (0x00000000000000000000000000009000) 
14'h0282 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000000000000; // D (0x00000000000000000000000000011000) 
14'h09eb : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100001000000000000; // D (0x00000000000000000000000000021000) 
14'h1f39 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000001000000000000; // D (0x00000000000000000000000000041000) 
14'h329d : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000001000000000000; // D (0x00000000000000000000000000081000) 
14'h2aa2 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000001000000000000; // D (0x00000000000000000000000000101000) 
14'h1adc : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000001000000000000; // D (0x00000000000000000000000000201000) 
14'h3957 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000001000000000000; // D (0x00000000000000000000000000401000) 
14'h3d36 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000001000000000000; // D (0x00000000000000000000000000801000) 
14'h35f4 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000001000000000000; // D (0x00000000000000000000000001001000) 
14'h2470 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000001000000000000; // D (0x00000000000000000000000002001000) 
14'h0778 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000001000000000000; // D (0x00000000000000000000000004001000) 
14'h021f : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000001000000000000; // D (0x00000000000000000000000008001000) 
14'h08d1 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001000000000000; // D (0x00000000000000000000000010001000) 
14'h1d4d : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000001000000000000; // D (0x00000000000000000000000020001000) 
14'h3675 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000001000000000000; // D (0x00000000000000000000000040001000) 
14'h2372 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000001000000000000; // D (0x00000000000000000000000080001000) 
14'h097c : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000001000000000000; // D (0x00000000000000000000000100001000) 
14'h1e17 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000001000000000000; // D (0x00000000000000000000000200001000) 
14'h30c1 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000001000000000000; // D (0x00000000000000000000000400001000) 
14'h2e1a : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000001000000000000; // D (0x00000000000000000000000800001000) 
14'h13ac : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000001000000000000; // D (0x00000000000000000000001000001000) 
14'h2bb7 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000001000000000000; // D (0x00000000000000000000002000001000) 
14'h18f6 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000001000000000000; // D (0x00000000000000000000004000001000) 
14'h3d03 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000001000000000000; // D (0x00000000000000000000008000001000) 
14'h359e : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000001000000000000; // D (0x00000000000000000000010000001000) 
14'h24a4 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000001000000000000; // D (0x00000000000000000000020000001000) 
14'h06d0 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000001000000000000; // D (0x00000000000000000000040000001000) 
14'h014f : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000001000000000000; // D (0x00000000000000000000080000001000) 
14'h0e71 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000001000000000000; // D (0x00000000000000000000100000001000) 
14'h100d : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000001000000000000; // D (0x00000000000000000000200000001000) 
14'h2cf5 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000001000000000000; // D (0x00000000000000000000400000001000) 
14'h1672 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000001000000000000; // D (0x00000000000000000000800000001000) 
14'h200b : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000001000000000000; // D (0x00000000000000000001000000001000) 
14'h0f8e : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000001000000000000; // D (0x00000000000000000002000000001000) 
14'h13f3 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000000; // D (0x00000000000000000004000000001000) 
14'h2b09 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000001000000000000; // D (0x00000000000000000008000000001000) 
14'h198a : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000001000000000000; // D (0x00000000000000000010000000001000) 
14'h3ffb : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000001000000000000; // D (0x00000000000000000020000000001000) 
14'h306e : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000001000000000000; // D (0x00000000000000000040000000001000) 
14'h2f44 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000001000000000000; // D (0x00000000000000000080000000001000) 
14'h1110 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000001000000000000; // D (0x00000000000000000100000000001000) 
14'h2ecf : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000001000000000000; // D (0x00000000000000000200000000001000) 
14'h1206 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000001000000000000; // D (0x00000000000000000400000000001000) 
14'h28e3 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000001000000000000; // D (0x00000000000000000800000000001000) 
14'h1e5e : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000001000000000000; // D (0x00000000000000001000000000001000) 
14'h3053 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000001000000000000; // D (0x00000000000000002000000000001000) 
14'h2f3e : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000001000000000000; // D (0x00000000000000004000000000001000) 
14'h11e4 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000001000000000000; // D (0x00000000000000008000000000001000) 
14'h2f27 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000001000000000000; // D (0x00000000000000010000000000001000) 
14'h11d6 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000001000000000000; // D (0x00000000000000020000000000001000) 
14'h2f43 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000001000000000000; // D (0x00000000000000040000000000001000) 
14'h111e : LOC =         127'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000001000000000000; // D (0x00000000000000080000000000001000) 
14'h2ed3 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000001000000000000; // D (0x00000000000000100000000000001000) 
14'h123e : LOC =         127'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000001000000000000; // D (0x00000000000000200000000000001000) 
14'h2893 : LOC =         127'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000001000000000000; // D (0x00000000000000400000000000001000) 
14'h1ebe : LOC =         127'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000001000000000000; // D (0x00000000000000800000000000001000) 
14'h3193 : LOC =         127'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000001000000000000; // D (0x00000000000001000000000000001000) 
14'h2cbe : LOC =         127'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000001000000000000; // D (0x00000000000002000000000000001000) 
14'h16e4 : LOC =         127'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000001000000000000; // D (0x00000000000004000000000000001000) 
14'h2127 : LOC =         127'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000001000000000000; // D (0x00000000000008000000000000001000) 
14'h0dd6 : LOC =         127'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000001000000000000; // D (0x00000000000010000000000000001000) 
14'h1743 : LOC =         127'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000001000000000000; // D (0x00000000000020000000000000001000) 
14'h2269 : LOC =         127'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000001000000000000; // D (0x00000000000040000000000000001000) 
14'h0b4a : LOC =         127'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000001000000000000; // D (0x00000000000080000000000000001000) 
14'h1a7b : LOC =         127'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000001000000000000; // D (0x00000000000100000000000000001000) 
14'h3819 : LOC =         127'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000001000000000000; // D (0x00000000000200000000000000001000) 
14'h3faa : LOC =         127'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000001000000000000; // D (0x00000000000400000000000000001000) 
14'h30cc : LOC =         127'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000001000000000000; // D (0x00000000000800000000000000001000) 
14'h2e00 : LOC =         127'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000001000000000000; // D (0x00000000001000000000000000001000) 
14'h1398 : LOC =         127'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000001000000000000; // D (0x00000000002000000000000000001000) 
14'h2bdf : LOC =         127'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000001000000000000; // D (0x00000000004000000000000000001000) 
14'h1826 : LOC =         127'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000001000000000000; // D (0x00000000008000000000000000001000) 
14'h3ca3 : LOC =         127'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000001000000000000; // D (0x00000000010000000000000000001000) 
14'h36de : LOC =         127'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000001000000000000; // D (0x00000000020000000000000000001000) 
14'h2224 : LOC =         127'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000; // D (0x00000000040000000000000000001000) 
14'h0bd0 : LOC =         127'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000; // D (0x00000000080000000000000000001000) 
14'h1b4f : LOC =         127'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000; // D (0x00000000100000000000000000001000) 
14'h3a71 : LOC =         127'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000; // D (0x00000000200000000000000000001000) 
14'h3b7a : LOC =         127'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000; // D (0x00000000400000000000000000001000) 
14'h396c : LOC =         127'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000; // D (0x00000000800000000000000000001000) 
14'h3d40 : LOC =         127'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000; // D (0x00000001000000000000000000001000) 
14'h3518 : LOC =         127'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000; // D (0x00000002000000000000000000001000) 
14'h25a8 : LOC =         127'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000; // D (0x00000004000000000000000000001000) 
14'h04c8 : LOC =         127'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000; // D (0x00000008000000000000000000001000) 
14'h057f : LOC =         127'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000; // D (0x00000010000000000000000000001000) 
14'h0611 : LOC =         127'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000; // D (0x00000020000000000000000000001000) 
14'h00cd : LOC =         127'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000; // D (0x00000040000000000000000000001000) 
14'h0d75 : LOC =         127'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000; // D (0x00000080000000000000000000001000) 
14'h1605 : LOC =         127'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000; // D (0x00000100000000000000000000001000) 
14'h20e5 : LOC =         127'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000; // D (0x00000200000000000000000000001000) 
14'h0e52 : LOC =         127'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000; // D (0x00000400000000000000000000001000) 
14'h104b : LOC =         127'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000; // D (0x00000800000000000000000000001000) 
14'h2c79 : LOC =         127'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000; // D (0x00001000000000000000000000001000) 
14'h176a : LOC =         127'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000; // D (0x00002000000000000000000000001000) 
14'h223b : LOC =         127'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000; // D (0x00004000000000000000000000001000) 
14'h0bee : LOC =         127'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000; // D (0x00008000000000000000000000001000) 
14'h1b33 : LOC =         127'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000; // D (0x00010000000000000000000000001000) 
14'h3a89 : LOC =         127'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000; // D (0x00020000000000000000000000001000) 
14'h3a8a : LOC =         127'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000; // D (0x00040000000000000000000000001000) 
14'h3a8c : LOC =         127'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000; // D (0x00080000000000000000000000001000) 
14'h3a80 : LOC =         127'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000; // D (0x00100000000000000000000000001000) 
14'h3a98 : LOC =         127'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000; // D (0x00200000000000000000000000001000) 
14'h3aa8 : LOC =         127'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000; // D (0x00400000000000000000000000001000) 
14'h3ac8 : LOC =         127'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000; // D (0x00800000000000000000000000001000) 
14'h3a08 : LOC =         127'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000; // D (0x01000000000000000000000000001000) 
14'h3b88 : LOC =         127'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000; // D (0x02000000000000000000000000001000) 
14'h3888 : LOC =         127'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000; // D (0x04000000000000000000000000001000) 
14'h3e88 : LOC =         127'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000; // D (0x08000000000000000000000000001000) 
14'h3288 : LOC =         127'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000; // D (0x10000000000000000000000000001000) 
14'h2a88 : LOC =         127'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000; // D (0x20000000000000000000000000001000) 
14'h1a88 : LOC =         127'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000; // D (0x40000000000000000000000000001000) 
14'h3667 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000; // S (0x00000000000000000000000000002000) 
14'h19de : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000; // D (0x00000000000000000000000000006000) 
14'h2a62 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000000000000; // D (0x0000000000000000000000000000a000) 
14'h0e6d : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000; // D (0x00000000000000000000000000012000) 
14'h0504 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010000000000000; // D (0x00000000000000000000000000022000) 
14'h13d6 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000010000000000000; // D (0x00000000000000000000000000042000) 
14'h3e72 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000010000000000000; // D (0x00000000000000000000000000082000) 
14'h264d : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000010000000000000; // D (0x00000000000000000000000000102000) 
14'h1633 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000010000000000000; // D (0x00000000000000000000000000202000) 
14'h35b8 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000010000000000000; // D (0x00000000000000000000000000402000) 
14'h31d9 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000010000000000000; // D (0x00000000000000000000000000802000) 
14'h391b : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000010000000000000; // D (0x00000000000000000000000001002000) 
14'h289f : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000010000000000000; // D (0x00000000000000000000000002002000) 
14'h0b97 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000010000000000000; // D (0x00000000000000000000000004002000) 
14'h0ef0 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000010000000000000; // D (0x00000000000000000000000008002000) 
14'h043e : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000010000000000000; // D (0x00000000000000000000000010002000) 
14'h11a2 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000010000000000000; // D (0x00000000000000000000000020002000) 
14'h3a9a : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000010000000000000; // D (0x00000000000000000000000040002000) 
14'h2f9d : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000010000000000000; // D (0x00000000000000000000000080002000) 
14'h0593 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000010000000000000; // D (0x00000000000000000000000100002000) 
14'h12f8 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000010000000000000; // D (0x00000000000000000000000200002000) 
14'h3c2e : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000010000000000000; // D (0x00000000000000000000000400002000) 
14'h22f5 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000010000000000000; // D (0x00000000000000000000000800002000) 
14'h1f43 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000010000000000000; // D (0x00000000000000000000001000002000) 
14'h2758 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000010000000000000; // D (0x00000000000000000000002000002000) 
14'h1419 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000010000000000000; // D (0x00000000000000000000004000002000) 
14'h31ec : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000010000000000000; // D (0x00000000000000000000008000002000) 
14'h3971 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000010000000000000; // D (0x00000000000000000000010000002000) 
14'h284b : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000010000000000000; // D (0x00000000000000000000020000002000) 
14'h0a3f : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000010000000000000; // D (0x00000000000000000000040000002000) 
14'h0da0 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000010000000000000; // D (0x00000000000000000000080000002000) 
14'h029e : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000010000000000000; // D (0x00000000000000000000100000002000) 
14'h1ce2 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000010000000000000; // D (0x00000000000000000000200000002000) 
14'h201a : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000010000000000000; // D (0x00000000000000000000400000002000) 
14'h1a9d : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000010000000000000; // D (0x00000000000000000000800000002000) 
14'h2ce4 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000010000000000000; // D (0x00000000000000000001000000002000) 
14'h0361 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000010000000000000; // D (0x00000000000000000002000000002000) 
14'h1f1c : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000010000000000000; // D (0x00000000000000000004000000002000) 
14'h27e6 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000010000000000000; // D (0x00000000000000000008000000002000) 
14'h1565 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000010000000000000; // D (0x00000000000000000010000000002000) 
14'h3314 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000010000000000000; // D (0x00000000000000000020000000002000) 
14'h3c81 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000010000000000000; // D (0x00000000000000000040000000002000) 
14'h23ab : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000010000000000000; // D (0x00000000000000000080000000002000) 
14'h1dff : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000010000000000000; // D (0x00000000000000000100000000002000) 
14'h2220 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000010000000000000; // D (0x00000000000000000200000000002000) 
14'h1ee9 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000010000000000000; // D (0x00000000000000000400000000002000) 
14'h240c : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000010000000000000; // D (0x00000000000000000800000000002000) 
14'h12b1 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000010000000000000; // D (0x00000000000000001000000000002000) 
14'h3cbc : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000010000000000000; // D (0x00000000000000002000000000002000) 
14'h23d1 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000010000000000000; // D (0x00000000000000004000000000002000) 
14'h1d0b : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000010000000000000; // D (0x00000000000000008000000000002000) 
14'h23c8 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000010000000000000; // D (0x00000000000000010000000000002000) 
14'h1d39 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000010000000000000; // D (0x00000000000000020000000000002000) 
14'h23ac : LOC =         127'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000010000000000000; // D (0x00000000000000040000000000002000) 
14'h1df1 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000010000000000000; // D (0x00000000000000080000000000002000) 
14'h223c : LOC =         127'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000010000000000000; // D (0x00000000000000100000000000002000) 
14'h1ed1 : LOC =         127'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000010000000000000; // D (0x00000000000000200000000000002000) 
14'h247c : LOC =         127'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000010000000000000; // D (0x00000000000000400000000000002000) 
14'h1251 : LOC =         127'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000010000000000000; // D (0x00000000000000800000000000002000) 
14'h3d7c : LOC =         127'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000010000000000000; // D (0x00000000000001000000000000002000) 
14'h2051 : LOC =         127'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000010000000000000; // D (0x00000000000002000000000000002000) 
14'h1a0b : LOC =         127'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000010000000000000; // D (0x00000000000004000000000000002000) 
14'h2dc8 : LOC =         127'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000010000000000000; // D (0x00000000000008000000000000002000) 
14'h0139 : LOC =         127'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000010000000000000; // D (0x00000000000010000000000000002000) 
14'h1bac : LOC =         127'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000010000000000000; // D (0x00000000000020000000000000002000) 
14'h2e86 : LOC =         127'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000010000000000000; // D (0x00000000000040000000000000002000) 
14'h07a5 : LOC =         127'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000010000000000000; // D (0x00000000000080000000000000002000) 
14'h1694 : LOC =         127'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000010000000000000; // D (0x00000000000100000000000000002000) 
14'h34f6 : LOC =         127'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000010000000000000; // D (0x00000000000200000000000000002000) 
14'h3345 : LOC =         127'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000010000000000000; // D (0x00000000000400000000000000002000) 
14'h3c23 : LOC =         127'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000010000000000000; // D (0x00000000000800000000000000002000) 
14'h22ef : LOC =         127'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000010000000000000; // D (0x00000000001000000000000000002000) 
14'h1f77 : LOC =         127'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000010000000000000; // D (0x00000000002000000000000000002000) 
14'h2730 : LOC =         127'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000010000000000000; // D (0x00000000004000000000000000002000) 
14'h14c9 : LOC =         127'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000010000000000000; // D (0x00000000008000000000000000002000) 
14'h304c : LOC =         127'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000010000000000000; // D (0x00000000010000000000000000002000) 
14'h3a31 : LOC =         127'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000010000000000000; // D (0x00000000020000000000000000002000) 
14'h2ecb : LOC =         127'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000; // D (0x00000000040000000000000000002000) 
14'h073f : LOC =         127'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000; // D (0x00000000080000000000000000002000) 
14'h17a0 : LOC =         127'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000; // D (0x00000000100000000000000000002000) 
14'h369e : LOC =         127'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000; // D (0x00000000200000000000000000002000) 
14'h3795 : LOC =         127'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000; // D (0x00000000400000000000000000002000) 
14'h3583 : LOC =         127'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000; // D (0x00000000800000000000000000002000) 
14'h31af : LOC =         127'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000; // D (0x00000001000000000000000000002000) 
14'h39f7 : LOC =         127'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000; // D (0x00000002000000000000000000002000) 
14'h2947 : LOC =         127'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000; // D (0x00000004000000000000000000002000) 
14'h0827 : LOC =         127'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000; // D (0x00000008000000000000000000002000) 
14'h0990 : LOC =         127'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000; // D (0x00000010000000000000000000002000) 
14'h0afe : LOC =         127'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000; // D (0x00000020000000000000000000002000) 
14'h0c22 : LOC =         127'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000; // D (0x00000040000000000000000000002000) 
14'h019a : LOC =         127'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000; // D (0x00000080000000000000000000002000) 
14'h1aea : LOC =         127'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000; // D (0x00000100000000000000000000002000) 
14'h2c0a : LOC =         127'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000; // D (0x00000200000000000000000000002000) 
14'h02bd : LOC =         127'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000; // D (0x00000400000000000000000000002000) 
14'h1ca4 : LOC =         127'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000; // D (0x00000800000000000000000000002000) 
14'h2096 : LOC =         127'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000; // D (0x00001000000000000000000000002000) 
14'h1b85 : LOC =         127'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000; // D (0x00002000000000000000000000002000) 
14'h2ed4 : LOC =         127'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000; // D (0x00004000000000000000000000002000) 
14'h0701 : LOC =         127'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000; // D (0x00008000000000000000000000002000) 
14'h17dc : LOC =         127'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000; // D (0x00010000000000000000000000002000) 
14'h3666 : LOC =         127'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000; // D (0x00020000000000000000000000002000) 
14'h3665 : LOC =         127'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000; // D (0x00040000000000000000000000002000) 
14'h3663 : LOC =         127'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000; // D (0x00080000000000000000000000002000) 
14'h366f : LOC =         127'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000; // D (0x00100000000000000000000000002000) 
14'h3677 : LOC =         127'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000; // D (0x00200000000000000000000000002000) 
14'h3647 : LOC =         127'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000; // D (0x00400000000000000000000000002000) 
14'h3627 : LOC =         127'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000; // D (0x00800000000000000000000000002000) 
14'h36e7 : LOC =         127'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000; // D (0x01000000000000000000000000002000) 
14'h3767 : LOC =         127'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000; // D (0x02000000000000000000000000002000) 
14'h3467 : LOC =         127'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000; // D (0x04000000000000000000000000002000) 
14'h3267 : LOC =         127'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000; // D (0x08000000000000000000000000002000) 
14'h3e67 : LOC =         127'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000; // D (0x10000000000000000000000000002000) 
14'h2667 : LOC =         127'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000; // D (0x20000000000000000000000000002000) 
14'h1667 : LOC =         127'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000; // D (0x40000000000000000000000000002000) 
14'h2fb9 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000; // S (0x00000000000000000000000000004000) 
14'h33bc : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000; // D (0x0000000000000000000000000000c000) 
14'h17b3 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000; // D (0x00000000000000000000000000014000) 
14'h1cda : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000; // D (0x00000000000000000000000000024000) 
14'h0a08 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000100000000000000; // D (0x00000000000000000000000000044000) 
14'h27ac : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000100000000000000; // D (0x00000000000000000000000000084000) 
14'h3f93 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000100000000000000; // D (0x00000000000000000000000000104000) 
14'h0fed : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000100000000000000; // D (0x00000000000000000000000000204000) 
14'h2c66 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000100000000000000; // D (0x00000000000000000000000000404000) 
14'h2807 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000100000000000000; // D (0x00000000000000000000000000804000) 
14'h20c5 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000100000000000000; // D (0x00000000000000000000000001004000) 
14'h3141 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000100000000000000; // D (0x00000000000000000000000002004000) 
14'h1249 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000100000000000000; // D (0x00000000000000000000000004004000) 
14'h172e : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000100000000000000; // D (0x00000000000000000000000008004000) 
14'h1de0 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000100000000000000; // D (0x00000000000000000000000010004000) 
14'h087c : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000100000000000000; // D (0x00000000000000000000000020004000) 
14'h2344 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000100000000000000; // D (0x00000000000000000000000040004000) 
14'h3643 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000100000000000000; // D (0x00000000000000000000000080004000) 
14'h1c4d : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000100000000000000; // D (0x00000000000000000000000100004000) 
14'h0b26 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000100000000000000; // D (0x00000000000000000000000200004000) 
14'h25f0 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000100000000000000; // D (0x00000000000000000000000400004000) 
14'h3b2b : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000100000000000000; // D (0x00000000000000000000000800004000) 
14'h069d : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000100000000000000; // D (0x00000000000000000000001000004000) 
14'h3e86 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000100000000000000; // D (0x00000000000000000000002000004000) 
14'h0dc7 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000100000000000000; // D (0x00000000000000000000004000004000) 
14'h2832 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000100000000000000; // D (0x00000000000000000000008000004000) 
14'h20af : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000100000000000000; // D (0x00000000000000000000010000004000) 
14'h3195 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000100000000000000; // D (0x00000000000000000000020000004000) 
14'h13e1 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000100000000000000; // D (0x00000000000000000000040000004000) 
14'h147e : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000100000000000000; // D (0x00000000000000000000080000004000) 
14'h1b40 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000100000000000000; // D (0x00000000000000000000100000004000) 
14'h053c : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000100000000000000; // D (0x00000000000000000000200000004000) 
14'h39c4 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000100000000000000; // D (0x00000000000000000000400000004000) 
14'h0343 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000100000000000000; // D (0x00000000000000000000800000004000) 
14'h353a : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000100000000000000; // D (0x00000000000000000001000000004000) 
14'h1abf : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000100000000000000; // D (0x00000000000000000002000000004000) 
14'h06c2 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000100000000000000; // D (0x00000000000000000004000000004000) 
14'h3e38 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000100000000000000; // D (0x00000000000000000008000000004000) 
14'h0cbb : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000100000000000000; // D (0x00000000000000000010000000004000) 
14'h2aca : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000100000000000000; // D (0x00000000000000000020000000004000) 
14'h255f : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000100000000000000; // D (0x00000000000000000040000000004000) 
14'h3a75 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000100000000000000; // D (0x00000000000000000080000000004000) 
14'h0421 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000100000000000000; // D (0x00000000000000000100000000004000) 
14'h3bfe : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000100000000000000; // D (0x00000000000000000200000000004000) 
14'h0737 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000100000000000000; // D (0x00000000000000000400000000004000) 
14'h3dd2 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000100000000000000; // D (0x00000000000000000800000000004000) 
14'h0b6f : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000100000000000000; // D (0x00000000000000001000000000004000) 
14'h2562 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000100000000000000; // D (0x00000000000000002000000000004000) 
14'h3a0f : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000100000000000000; // D (0x00000000000000004000000000004000) 
14'h04d5 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000100000000000000; // D (0x00000000000000008000000000004000) 
14'h3a16 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000100000000000000; // D (0x00000000000000010000000000004000) 
14'h04e7 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000100000000000000; // D (0x00000000000000020000000000004000) 
14'h3a72 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000100000000000000; // D (0x00000000000000040000000000004000) 
14'h042f : LOC =         127'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000100000000000000; // D (0x00000000000000080000000000004000) 
14'h3be2 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000100000000000000; // D (0x00000000000000100000000000004000) 
14'h070f : LOC =         127'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000100000000000000; // D (0x00000000000000200000000000004000) 
14'h3da2 : LOC =         127'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000100000000000000; // D (0x00000000000000400000000000004000) 
14'h0b8f : LOC =         127'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000100000000000000; // D (0x00000000000000800000000000004000) 
14'h24a2 : LOC =         127'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000100000000000000; // D (0x00000000000001000000000000004000) 
14'h398f : LOC =         127'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000100000000000000; // D (0x00000000000002000000000000004000) 
14'h03d5 : LOC =         127'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000100000000000000; // D (0x00000000000004000000000000004000) 
14'h3416 : LOC =         127'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000100000000000000; // D (0x00000000000008000000000000004000) 
14'h18e7 : LOC =         127'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000100000000000000; // D (0x00000000000010000000000000004000) 
14'h0272 : LOC =         127'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000100000000000000; // D (0x00000000000020000000000000004000) 
14'h3758 : LOC =         127'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000100000000000000; // D (0x00000000000040000000000000004000) 
14'h1e7b : LOC =         127'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000100000000000000; // D (0x00000000000080000000000000004000) 
14'h0f4a : LOC =         127'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000100000000000000; // D (0x00000000000100000000000000004000) 
14'h2d28 : LOC =         127'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000100000000000000; // D (0x00000000000200000000000000004000) 
14'h2a9b : LOC =         127'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000100000000000000; // D (0x00000000000400000000000000004000) 
14'h25fd : LOC =         127'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000100000000000000; // D (0x00000000000800000000000000004000) 
14'h3b31 : LOC =         127'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000100000000000000; // D (0x00000000001000000000000000004000) 
14'h06a9 : LOC =         127'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000100000000000000; // D (0x00000000002000000000000000004000) 
14'h3eee : LOC =         127'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000100000000000000; // D (0x00000000004000000000000000004000) 
14'h0d17 : LOC =         127'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000100000000000000; // D (0x00000000008000000000000000004000) 
14'h2992 : LOC =         127'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000100000000000000; // D (0x00000000010000000000000000004000) 
14'h23ef : LOC =         127'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000100000000000000; // D (0x00000000020000000000000000004000) 
14'h3715 : LOC =         127'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000; // D (0x00000000040000000000000000004000) 
14'h1ee1 : LOC =         127'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000; // D (0x00000000080000000000000000004000) 
14'h0e7e : LOC =         127'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000; // D (0x00000000100000000000000000004000) 
14'h2f40 : LOC =         127'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000; // D (0x00000000200000000000000000004000) 
14'h2e4b : LOC =         127'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000; // D (0x00000000400000000000000000004000) 
14'h2c5d : LOC =         127'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000; // D (0x00000000800000000000000000004000) 
14'h2871 : LOC =         127'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000; // D (0x00000001000000000000000000004000) 
14'h2029 : LOC =         127'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000; // D (0x00000002000000000000000000004000) 
14'h3099 : LOC =         127'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000; // D (0x00000004000000000000000000004000) 
14'h11f9 : LOC =         127'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000; // D (0x00000008000000000000000000004000) 
14'h104e : LOC =         127'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000; // D (0x00000010000000000000000000004000) 
14'h1320 : LOC =         127'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000; // D (0x00000020000000000000000000004000) 
14'h15fc : LOC =         127'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000; // D (0x00000040000000000000000000004000) 
14'h1844 : LOC =         127'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000; // D (0x00000080000000000000000000004000) 
14'h0334 : LOC =         127'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000; // D (0x00000100000000000000000000004000) 
14'h35d4 : LOC =         127'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000; // D (0x00000200000000000000000000004000) 
14'h1b63 : LOC =         127'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000; // D (0x00000400000000000000000000004000) 
14'h057a : LOC =         127'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000; // D (0x00000800000000000000000000004000) 
14'h3948 : LOC =         127'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000; // D (0x00001000000000000000000000004000) 
14'h025b : LOC =         127'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000; // D (0x00002000000000000000000000004000) 
14'h370a : LOC =         127'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000; // D (0x00004000000000000000000000004000) 
14'h1edf : LOC =         127'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000; // D (0x00008000000000000000000000004000) 
14'h0e02 : LOC =         127'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000; // D (0x00010000000000000000000000004000) 
14'h2fb8 : LOC =         127'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000; // D (0x00020000000000000000000000004000) 
14'h2fbb : LOC =         127'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000; // D (0x00040000000000000000000000004000) 
14'h2fbd : LOC =         127'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000; // D (0x00080000000000000000000000004000) 
14'h2fb1 : LOC =         127'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000; // D (0x00100000000000000000000000004000) 
14'h2fa9 : LOC =         127'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000; // D (0x00200000000000000000000000004000) 
14'h2f99 : LOC =         127'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000; // D (0x00400000000000000000000000004000) 
14'h2ff9 : LOC =         127'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000; // D (0x00800000000000000000000000004000) 
14'h2f39 : LOC =         127'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000; // D (0x01000000000000000000000000004000) 
14'h2eb9 : LOC =         127'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000; // D (0x02000000000000000000000000004000) 
14'h2db9 : LOC =         127'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000; // D (0x04000000000000000000000000004000) 
14'h2bb9 : LOC =         127'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000; // D (0x08000000000000000000000000004000) 
14'h27b9 : LOC =         127'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000; // D (0x10000000000000000000000000004000) 
14'h3fb9 : LOC =         127'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000; // D (0x20000000000000000000000000004000) 
14'h0fb9 : LOC =         127'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000; // D (0x40000000000000000000000000004000) 
14'h1c05 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000; // S (0x00000000000000000000000000008000) 
14'h240f : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000; // D (0x00000000000000000000000000018000) 
14'h2f66 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000000000000000; // D (0x00000000000000000000000000028000) 
14'h39b4 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000; // D (0x00000000000000000000000000048000) 
14'h1410 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000000000000000; // D (0x00000000000000000000000000088000) 
14'h0c2f : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100001000000000000000; // D (0x00000000000000000000000000108000) 
14'h3c51 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000001000000000000000; // D (0x00000000000000000000000000208000) 
14'h1fda : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000001000000000000000; // D (0x00000000000000000000000000408000) 
14'h1bbb : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000001000000000000000; // D (0x00000000000000000000000000808000) 
14'h1379 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000001000000000000000; // D (0x00000000000000000000000001008000) 
14'h02fd : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000001000000000000000; // D (0x00000000000000000000000002008000) 
14'h21f5 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000001000000000000000; // D (0x00000000000000000000000004008000) 
14'h2492 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000001000000000000000; // D (0x00000000000000000000000008008000) 
14'h2e5c : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000001000000000000000; // D (0x00000000000000000000000010008000) 
14'h3bc0 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000001000000000000000; // D (0x00000000000000000000000020008000) 
14'h10f8 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000001000000000000000; // D (0x00000000000000000000000040008000) 
14'h05ff : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001000000000000000; // D (0x00000000000000000000000080008000) 
14'h2ff1 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000001000000000000000; // D (0x00000000000000000000000100008000) 
14'h389a : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000001000000000000000; // D (0x00000000000000000000000200008000) 
14'h164c : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000001000000000000000; // D (0x00000000000000000000000400008000) 
14'h0897 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000001000000000000000; // D (0x00000000000000000000000800008000) 
14'h3521 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000001000000000000000; // D (0x00000000000000000000001000008000) 
14'h0d3a : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000001000000000000000; // D (0x00000000000000000000002000008000) 
14'h3e7b : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000001000000000000000; // D (0x00000000000000000000004000008000) 
14'h1b8e : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000001000000000000000; // D (0x00000000000000000000008000008000) 
14'h1313 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000001000000000000000; // D (0x00000000000000000000010000008000) 
14'h0229 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000001000000000000000; // D (0x00000000000000000000020000008000) 
14'h205d : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000001000000000000000; // D (0x00000000000000000000040000008000) 
14'h27c2 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000001000000000000000; // D (0x00000000000000000000080000008000) 
14'h28fc : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000001000000000000000; // D (0x00000000000000000000100000008000) 
14'h3680 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000001000000000000000; // D (0x00000000000000000000200000008000) 
14'h0a78 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000001000000000000000; // D (0x00000000000000000000400000008000) 
14'h30ff : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000001000000000000000; // D (0x00000000000000000000800000008000) 
14'h0686 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000001000000000000000; // D (0x00000000000000000001000000008000) 
14'h2903 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000001000000000000000; // D (0x00000000000000000002000000008000) 
14'h357e : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000001000000000000000; // D (0x00000000000000000004000000008000) 
14'h0d84 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000001000000000000000; // D (0x00000000000000000008000000008000) 
14'h3f07 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000001000000000000000; // D (0x00000000000000000010000000008000) 
14'h1976 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000000000; // D (0x00000000000000000020000000008000) 
14'h16e3 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000001000000000000000; // D (0x00000000000000000040000000008000) 
14'h09c9 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000001000000000000000; // D (0x00000000000000000080000000008000) 
14'h379d : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000001000000000000000; // D (0x00000000000000000100000000008000) 
14'h0842 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000001000000000000000; // D (0x00000000000000000200000000008000) 
14'h348b : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000001000000000000000; // D (0x00000000000000000400000000008000) 
14'h0e6e : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000001000000000000000; // D (0x00000000000000000800000000008000) 
14'h38d3 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000001000000000000000; // D (0x00000000000000001000000000008000) 
14'h16de : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000001000000000000000; // D (0x00000000000000002000000000008000) 
14'h09b3 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000001000000000000000; // D (0x00000000000000004000000000008000) 
14'h3769 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000001000000000000000; // D (0x00000000000000008000000000008000) 
14'h09aa : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000001000000000000000; // D (0x00000000000000010000000000008000) 
14'h375b : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000001000000000000000; // D (0x00000000000000020000000000008000) 
14'h09ce : LOC =         127'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000001000000000000000; // D (0x00000000000000040000000000008000) 
14'h3793 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000001000000000000000; // D (0x00000000000000080000000000008000) 
14'h085e : LOC =         127'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000001000000000000000; // D (0x00000000000000100000000000008000) 
14'h34b3 : LOC =         127'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000001000000000000000; // D (0x00000000000000200000000000008000) 
14'h0e1e : LOC =         127'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000001000000000000000; // D (0x00000000000000400000000000008000) 
14'h3833 : LOC =         127'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000001000000000000000; // D (0x00000000000000800000000000008000) 
14'h171e : LOC =         127'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000001000000000000000; // D (0x00000000000001000000000000008000) 
14'h0a33 : LOC =         127'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000001000000000000000; // D (0x00000000000002000000000000008000) 
14'h3069 : LOC =         127'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000001000000000000000; // D (0x00000000000004000000000000008000) 
14'h07aa : LOC =         127'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000001000000000000000; // D (0x00000000000008000000000000008000) 
14'h2b5b : LOC =         127'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000001000000000000000; // D (0x00000000000010000000000000008000) 
14'h31ce : LOC =         127'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000001000000000000000; // D (0x00000000000020000000000000008000) 
14'h04e4 : LOC =         127'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000001000000000000000; // D (0x00000000000040000000000000008000) 
14'h2dc7 : LOC =         127'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000001000000000000000; // D (0x00000000000080000000000000008000) 
14'h3cf6 : LOC =         127'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000001000000000000000; // D (0x00000000000100000000000000008000) 
14'h1e94 : LOC =         127'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000001000000000000000; // D (0x00000000000200000000000000008000) 
14'h1927 : LOC =         127'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000001000000000000000; // D (0x00000000000400000000000000008000) 
14'h1641 : LOC =         127'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000001000000000000000; // D (0x00000000000800000000000000008000) 
14'h088d : LOC =         127'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000001000000000000000; // D (0x00000000001000000000000000008000) 
14'h3515 : LOC =         127'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000001000000000000000; // D (0x00000000002000000000000000008000) 
14'h0d52 : LOC =         127'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000001000000000000000; // D (0x00000000004000000000000000008000) 
14'h3eab : LOC =         127'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000001000000000000000; // D (0x00000000008000000000000000008000) 
14'h1a2e : LOC =         127'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000001000000000000000; // D (0x00000000010000000000000000008000) 
14'h1053 : LOC =         127'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000001000000000000000; // D (0x00000000020000000000000000008000) 
14'h04a9 : LOC =         127'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000; // D (0x00000000040000000000000000008000) 
14'h2d5d : LOC =         127'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000; // D (0x00000000080000000000000000008000) 
14'h3dc2 : LOC =         127'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000; // D (0x00000000100000000000000000008000) 
14'h1cfc : LOC =         127'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000; // D (0x00000000200000000000000000008000) 
14'h1df7 : LOC =         127'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000; // D (0x00000000400000000000000000008000) 
14'h1fe1 : LOC =         127'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000; // D (0x00000000800000000000000000008000) 
14'h1bcd : LOC =         127'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000; // D (0x00000001000000000000000000008000) 
14'h1395 : LOC =         127'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000; // D (0x00000002000000000000000000008000) 
14'h0325 : LOC =         127'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000; // D (0x00000004000000000000000000008000) 
14'h2245 : LOC =         127'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000; // D (0x00000008000000000000000000008000) 
14'h23f2 : LOC =         127'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000; // D (0x00000010000000000000000000008000) 
14'h209c : LOC =         127'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000; // D (0x00000020000000000000000000008000) 
14'h2640 : LOC =         127'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000; // D (0x00000040000000000000000000008000) 
14'h2bf8 : LOC =         127'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000; // D (0x00000080000000000000000000008000) 
14'h3088 : LOC =         127'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000; // D (0x00000100000000000000000000008000) 
14'h0668 : LOC =         127'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000; // D (0x00000200000000000000000000008000) 
14'h28df : LOC =         127'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000; // D (0x00000400000000000000000000008000) 
14'h36c6 : LOC =         127'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000; // D (0x00000800000000000000000000008000) 
14'h0af4 : LOC =         127'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000; // D (0x00001000000000000000000000008000) 
14'h31e7 : LOC =         127'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000; // D (0x00002000000000000000000000008000) 
14'h04b6 : LOC =         127'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000; // D (0x00004000000000000000000000008000) 
14'h2d63 : LOC =         127'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000; // D (0x00008000000000000000000000008000) 
14'h3dbe : LOC =         127'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000; // D (0x00010000000000000000000000008000) 
14'h1c04 : LOC =         127'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000; // D (0x00020000000000000000000000008000) 
14'h1c07 : LOC =         127'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000; // D (0x00040000000000000000000000008000) 
14'h1c01 : LOC =         127'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000; // D (0x00080000000000000000000000008000) 
14'h1c0d : LOC =         127'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000; // D (0x00100000000000000000000000008000) 
14'h1c15 : LOC =         127'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000; // D (0x00200000000000000000000000008000) 
14'h1c25 : LOC =         127'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000; // D (0x00400000000000000000000000008000) 
14'h1c45 : LOC =         127'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000; // D (0x00800000000000000000000000008000) 
14'h1c85 : LOC =         127'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000; // D (0x01000000000000000000000000008000) 
14'h1d05 : LOC =         127'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000; // D (0x02000000000000000000000000008000) 
14'h1e05 : LOC =         127'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000; // D (0x04000000000000000000000000008000) 
14'h1805 : LOC =         127'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000; // D (0x08000000000000000000000000008000) 
14'h1405 : LOC =         127'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000; // D (0x10000000000000000000000000008000) 
14'h0c05 : LOC =         127'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000; // D (0x20000000000000000000000000008000) 
14'h3c05 : LOC =         127'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000; // D (0x40000000000000000000000000008000) 
14'h380a : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000; // S (0x00000000000000000000000000010000) 
14'h0b69 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000; // D (0x00000000000000000000000000030000) 
14'h1dbb : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000000000000000; // D (0x00000000000000000000000000050000) 
14'h301f : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000; // D (0x00000000000000000000000000090000) 
14'h2820 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010000000000000000; // D (0x00000000000000000000000000110000) 
14'h185e : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000010000000000000000; // D (0x00000000000000000000000000210000) 
14'h3bd5 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000010000000000000000; // D (0x00000000000000000000000000410000) 
14'h3fb4 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000010000000000000000; // D (0x00000000000000000000000000810000) 
14'h3776 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000010000000000000000; // D (0x00000000000000000000000001010000) 
14'h26f2 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000010000000000000000; // D (0x00000000000000000000000002010000) 
14'h05fa : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000010000000000000000; // D (0x00000000000000000000000004010000) 
14'h009d : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000010000000000000000; // D (0x00000000000000000000000008010000) 
14'h0a53 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000010000000000000000; // D (0x00000000000000000000000010010000) 
14'h1fcf : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000010000000000000000; // D (0x00000000000000000000000020010000) 
14'h34f7 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000010000000000000000; // D (0x00000000000000000000000040010000) 
14'h21f0 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000010000000000000000; // D (0x00000000000000000000000080010000) 
14'h0bfe : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000010000000000000000; // D (0x00000000000000000000000100010000) 
14'h1c95 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000010000000000000000; // D (0x00000000000000000000000200010000) 
14'h3243 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000010000000000000000; // D (0x00000000000000000000000400010000) 
14'h2c98 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000010000000000000000; // D (0x00000000000000000000000800010000) 
14'h112e : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000010000000000000000; // D (0x00000000000000000000001000010000) 
14'h2935 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000010000000000000000; // D (0x00000000000000000000002000010000) 
14'h1a74 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000010000000000000000; // D (0x00000000000000000000004000010000) 
14'h3f81 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000010000000000000000; // D (0x00000000000000000000008000010000) 
14'h371c : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000010000000000000000; // D (0x00000000000000000000010000010000) 
14'h2626 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000010000000000000000; // D (0x00000000000000000000020000010000) 
14'h0452 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000010000000000000000; // D (0x00000000000000000000040000010000) 
14'h03cd : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000010000000000000000; // D (0x00000000000000000000080000010000) 
14'h0cf3 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000010000000000000000; // D (0x00000000000000000000100000010000) 
14'h128f : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000010000000000000000; // D (0x00000000000000000000200000010000) 
14'h2e77 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000010000000000000000; // D (0x00000000000000000000400000010000) 
14'h14f0 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000010000000000000000; // D (0x00000000000000000000800000010000) 
14'h2289 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000010000000000000000; // D (0x00000000000000000001000000010000) 
14'h0d0c : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000010000000000000000; // D (0x00000000000000000002000000010000) 
14'h1171 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000010000000000000000; // D (0x00000000000000000004000000010000) 
14'h298b : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000010000000000000000; // D (0x00000000000000000008000000010000) 
14'h1b08 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000010000000000000000; // D (0x00000000000000000010000000010000) 
14'h3d79 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000010000000000000000; // D (0x00000000000000000020000000010000) 
14'h32ec : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000010000000000000000; // D (0x00000000000000000040000000010000) 
14'h2dc6 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000010000000000000000; // D (0x00000000000000000080000000010000) 
14'h1392 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000010000000000000000; // D (0x00000000000000000100000000010000) 
14'h2c4d : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000010000000000000000; // D (0x00000000000000000200000000010000) 
14'h1084 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000010000000000000000; // D (0x00000000000000000400000000010000) 
14'h2a61 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000010000000000000000; // D (0x00000000000000000800000000010000) 
14'h1cdc : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000010000000000000000; // D (0x00000000000000001000000000010000) 
14'h32d1 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000010000000000000000; // D (0x00000000000000002000000000010000) 
14'h2dbc : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000010000000000000000; // D (0x00000000000000004000000000010000) 
14'h1366 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000010000000000000000; // D (0x00000000000000008000000000010000) 
14'h2da5 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000010000000000000000; // D (0x00000000000000010000000000010000) 
14'h1354 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000010000000000000000; // D (0x00000000000000020000000000010000) 
14'h2dc1 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000010000000000000000; // D (0x00000000000000040000000000010000) 
14'h139c : LOC =         127'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000010000000000000000; // D (0x00000000000000080000000000010000) 
14'h2c51 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000010000000000000000; // D (0x00000000000000100000000000010000) 
14'h10bc : LOC =         127'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000010000000000000000; // D (0x00000000000000200000000000010000) 
14'h2a11 : LOC =         127'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000010000000000000000; // D (0x00000000000000400000000000010000) 
14'h1c3c : LOC =         127'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000010000000000000000; // D (0x00000000000000800000000000010000) 
14'h3311 : LOC =         127'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000010000000000000000; // D (0x00000000000001000000000000010000) 
14'h2e3c : LOC =         127'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000010000000000000000; // D (0x00000000000002000000000000010000) 
14'h1466 : LOC =         127'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000010000000000000000; // D (0x00000000000004000000000000010000) 
14'h23a5 : LOC =         127'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000010000000000000000; // D (0x00000000000008000000000000010000) 
14'h0f54 : LOC =         127'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000010000000000000000; // D (0x00000000000010000000000000010000) 
14'h15c1 : LOC =         127'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000010000000000000000; // D (0x00000000000020000000000000010000) 
14'h20eb : LOC =         127'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000010000000000000000; // D (0x00000000000040000000000000010000) 
14'h09c8 : LOC =         127'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000010000000000000000; // D (0x00000000000080000000000000010000) 
14'h18f9 : LOC =         127'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000010000000000000000; // D (0x00000000000100000000000000010000) 
14'h3a9b : LOC =         127'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000010000000000000000; // D (0x00000000000200000000000000010000) 
14'h3d28 : LOC =         127'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000010000000000000000; // D (0x00000000000400000000000000010000) 
14'h324e : LOC =         127'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000010000000000000000; // D (0x00000000000800000000000000010000) 
14'h2c82 : LOC =         127'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000010000000000000000; // D (0x00000000001000000000000000010000) 
14'h111a : LOC =         127'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000010000000000000000; // D (0x00000000002000000000000000010000) 
14'h295d : LOC =         127'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000010000000000000000; // D (0x00000000004000000000000000010000) 
14'h1aa4 : LOC =         127'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000010000000000000000; // D (0x00000000008000000000000000010000) 
14'h3e21 : LOC =         127'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000010000000000000000; // D (0x00000000010000000000000000010000) 
14'h345c : LOC =         127'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000010000000000000000; // D (0x00000000020000000000000000010000) 
14'h20a6 : LOC =         127'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000; // D (0x00000000040000000000000000010000) 
14'h0952 : LOC =         127'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000; // D (0x00000000080000000000000000010000) 
14'h19cd : LOC =         127'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000; // D (0x00000000100000000000000000010000) 
14'h38f3 : LOC =         127'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000; // D (0x00000000200000000000000000010000) 
14'h39f8 : LOC =         127'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000; // D (0x00000000400000000000000000010000) 
14'h3bee : LOC =         127'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000; // D (0x00000000800000000000000000010000) 
14'h3fc2 : LOC =         127'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000; // D (0x00000001000000000000000000010000) 
14'h379a : LOC =         127'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000; // D (0x00000002000000000000000000010000) 
14'h272a : LOC =         127'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000; // D (0x00000004000000000000000000010000) 
14'h064a : LOC =         127'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000; // D (0x00000008000000000000000000010000) 
14'h07fd : LOC =         127'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000; // D (0x00000010000000000000000000010000) 
14'h0493 : LOC =         127'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000; // D (0x00000020000000000000000000010000) 
14'h024f : LOC =         127'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000; // D (0x00000040000000000000000000010000) 
14'h0ff7 : LOC =         127'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000; // D (0x00000080000000000000000000010000) 
14'h1487 : LOC =         127'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000; // D (0x00000100000000000000000000010000) 
14'h2267 : LOC =         127'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000; // D (0x00000200000000000000000000010000) 
14'h0cd0 : LOC =         127'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000; // D (0x00000400000000000000000000010000) 
14'h12c9 : LOC =         127'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000; // D (0x00000800000000000000000000010000) 
14'h2efb : LOC =         127'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000; // D (0x00001000000000000000000000010000) 
14'h15e8 : LOC =         127'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000; // D (0x00002000000000000000000000010000) 
14'h20b9 : LOC =         127'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000; // D (0x00004000000000000000000000010000) 
14'h096c : LOC =         127'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000; // D (0x00008000000000000000000000010000) 
14'h19b1 : LOC =         127'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000; // D (0x00010000000000000000000000010000) 
14'h380b : LOC =         127'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000; // D (0x00020000000000000000000000010000) 
14'h3808 : LOC =         127'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000; // D (0x00040000000000000000000000010000) 
14'h380e : LOC =         127'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000; // D (0x00080000000000000000000000010000) 
14'h3802 : LOC =         127'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000; // D (0x00100000000000000000000000010000) 
14'h381a : LOC =         127'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000; // D (0x00200000000000000000000000010000) 
14'h382a : LOC =         127'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000; // D (0x00400000000000000000000000010000) 
14'h384a : LOC =         127'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000; // D (0x00800000000000000000000000010000) 
14'h388a : LOC =         127'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000; // D (0x01000000000000000000000000010000) 
14'h390a : LOC =         127'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000; // D (0x02000000000000000000000000010000) 
14'h3a0a : LOC =         127'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000; // D (0x04000000000000000000000000010000) 
14'h3c0a : LOC =         127'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000; // D (0x08000000000000000000000000010000) 
14'h300a : LOC =         127'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000; // D (0x10000000000000000000000000010000) 
14'h280a : LOC =         127'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000; // D (0x20000000000000000000000000010000) 
14'h180a : LOC =         127'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000; // D (0x40000000000000000000000000010000) 
14'h3363 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000; // S (0x00000000000000000000000000020000) 
14'h16d2 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000; // D (0x00000000000000000000000000060000) 
14'h3b76 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000; // D (0x000000000000000000000000000a0000) 
14'h2349 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000; // D (0x00000000000000000000000000120000) 
14'h1337 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000100000000000000000; // D (0x00000000000000000000000000220000) 
14'h30bc : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000100000000000000000; // D (0x00000000000000000000000000420000) 
14'h34dd : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000100000000000000000; // D (0x00000000000000000000000000820000) 
14'h3c1f : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000100000000000000000; // D (0x00000000000000000000000001020000) 
14'h2d9b : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000100000000000000000; // D (0x00000000000000000000000002020000) 
14'h0e93 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000100000000000000000; // D (0x00000000000000000000000004020000) 
14'h0bf4 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000100000000000000000; // D (0x00000000000000000000000008020000) 
14'h013a : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000100000000000000000; // D (0x00000000000000000000000010020000) 
14'h14a6 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000100000000000000000; // D (0x00000000000000000000000020020000) 
14'h3f9e : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000100000000000000000; // D (0x00000000000000000000000040020000) 
14'h2a99 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000100000000000000000; // D (0x00000000000000000000000080020000) 
14'h0097 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000100000000000000000; // D (0x00000000000000000000000100020000) 
14'h17fc : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000100000000000000000; // D (0x00000000000000000000000200020000) 
14'h392a : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000100000000000000000; // D (0x00000000000000000000000400020000) 
14'h27f1 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000100000000000000000; // D (0x00000000000000000000000800020000) 
14'h1a47 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000100000000000000000; // D (0x00000000000000000000001000020000) 
14'h225c : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000100000000000000000; // D (0x00000000000000000000002000020000) 
14'h111d : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000100000000000000000; // D (0x00000000000000000000004000020000) 
14'h34e8 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000100000000000000000; // D (0x00000000000000000000008000020000) 
14'h3c75 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000100000000000000000; // D (0x00000000000000000000010000020000) 
14'h2d4f : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000100000000000000000; // D (0x00000000000000000000020000020000) 
14'h0f3b : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000100000000000000000; // D (0x00000000000000000000040000020000) 
14'h08a4 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000100000000000000000; // D (0x00000000000000000000080000020000) 
14'h079a : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000100000000000000000; // D (0x00000000000000000000100000020000) 
14'h19e6 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000100000000000000000; // D (0x00000000000000000000200000020000) 
14'h251e : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000100000000000000000; // D (0x00000000000000000000400000020000) 
14'h1f99 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000100000000000000000; // D (0x00000000000000000000800000020000) 
14'h29e0 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000100000000000000000; // D (0x00000000000000000001000000020000) 
14'h0665 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000100000000000000000; // D (0x00000000000000000002000000020000) 
14'h1a18 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000100000000000000000; // D (0x00000000000000000004000000020000) 
14'h22e2 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000100000000000000000; // D (0x00000000000000000008000000020000) 
14'h1061 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000100000000000000000; // D (0x00000000000000000010000000020000) 
14'h3610 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000100000000000000000; // D (0x00000000000000000020000000020000) 
14'h3985 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000100000000000000000; // D (0x00000000000000000040000000020000) 
14'h26af : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000100000000000000000; // D (0x00000000000000000080000000020000) 
14'h18fb : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000100000000000000000; // D (0x00000000000000000100000000020000) 
14'h2724 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000100000000000000000; // D (0x00000000000000000200000000020000) 
14'h1bed : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000100000000000000000; // D (0x00000000000000000400000000020000) 
14'h2108 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000100000000000000000; // D (0x00000000000000000800000000020000) 
14'h17b5 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000100000000000000000; // D (0x00000000000000001000000000020000) 
14'h39b8 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000100000000000000000; // D (0x00000000000000002000000000020000) 
14'h26d5 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000100000000000000000; // D (0x00000000000000004000000000020000) 
14'h180f : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000100000000000000000; // D (0x00000000000000008000000000020000) 
14'h26cc : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000100000000000000000; // D (0x00000000000000010000000000020000) 
14'h183d : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000100000000000000000; // D (0x00000000000000020000000000020000) 
14'h26a8 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000100000000000000000; // D (0x00000000000000040000000000020000) 
14'h18f5 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000100000000000000000; // D (0x00000000000000080000000000020000) 
14'h2738 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000100000000000000000; // D (0x00000000000000100000000000020000) 
14'h1bd5 : LOC =         127'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000100000000000000000; // D (0x00000000000000200000000000020000) 
14'h2178 : LOC =         127'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000100000000000000000; // D (0x00000000000000400000000000020000) 
14'h1755 : LOC =         127'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000100000000000000000; // D (0x00000000000000800000000000020000) 
14'h3878 : LOC =         127'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000100000000000000000; // D (0x00000000000001000000000000020000) 
14'h2555 : LOC =         127'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000100000000000000000; // D (0x00000000000002000000000000020000) 
14'h1f0f : LOC =         127'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000100000000000000000; // D (0x00000000000004000000000000020000) 
14'h28cc : LOC =         127'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000100000000000000000; // D (0x00000000000008000000000000020000) 
14'h043d : LOC =         127'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000100000000000000000; // D (0x00000000000010000000000000020000) 
14'h1ea8 : LOC =         127'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000100000000000000000; // D (0x00000000000020000000000000020000) 
14'h2b82 : LOC =         127'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000100000000000000000; // D (0x00000000000040000000000000020000) 
14'h02a1 : LOC =         127'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000100000000000000000; // D (0x00000000000080000000000000020000) 
14'h1390 : LOC =         127'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000100000000000000000; // D (0x00000000000100000000000000020000) 
14'h31f2 : LOC =         127'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000100000000000000000; // D (0x00000000000200000000000000020000) 
14'h3641 : LOC =         127'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000100000000000000000; // D (0x00000000000400000000000000020000) 
14'h3927 : LOC =         127'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000100000000000000000; // D (0x00000000000800000000000000020000) 
14'h27eb : LOC =         127'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000100000000000000000; // D (0x00000000001000000000000000020000) 
14'h1a73 : LOC =         127'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000100000000000000000; // D (0x00000000002000000000000000020000) 
14'h2234 : LOC =         127'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000100000000000000000; // D (0x00000000004000000000000000020000) 
14'h11cd : LOC =         127'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000100000000000000000; // D (0x00000000008000000000000000020000) 
14'h3548 : LOC =         127'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000100000000000000000; // D (0x00000000010000000000000000020000) 
14'h3f35 : LOC =         127'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000100000000000000000; // D (0x00000000020000000000000000020000) 
14'h2bcf : LOC =         127'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000; // D (0x00000000040000000000000000020000) 
14'h023b : LOC =         127'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000; // D (0x00000000080000000000000000020000) 
14'h12a4 : LOC =         127'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000; // D (0x00000000100000000000000000020000) 
14'h339a : LOC =         127'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000; // D (0x00000000200000000000000000020000) 
14'h3291 : LOC =         127'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000; // D (0x00000000400000000000000000020000) 
14'h3087 : LOC =         127'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000; // D (0x00000000800000000000000000020000) 
14'h34ab : LOC =         127'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000; // D (0x00000001000000000000000000020000) 
14'h3cf3 : LOC =         127'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000; // D (0x00000002000000000000000000020000) 
14'h2c43 : LOC =         127'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000; // D (0x00000004000000000000000000020000) 
14'h0d23 : LOC =         127'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000; // D (0x00000008000000000000000000020000) 
14'h0c94 : LOC =         127'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000; // D (0x00000010000000000000000000020000) 
14'h0ffa : LOC =         127'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000; // D (0x00000020000000000000000000020000) 
14'h0926 : LOC =         127'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000; // D (0x00000040000000000000000000020000) 
14'h049e : LOC =         127'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000; // D (0x00000080000000000000000000020000) 
14'h1fee : LOC =         127'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000; // D (0x00000100000000000000000000020000) 
14'h290e : LOC =         127'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000; // D (0x00000200000000000000000000020000) 
14'h07b9 : LOC =         127'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000; // D (0x00000400000000000000000000020000) 
14'h19a0 : LOC =         127'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000; // D (0x00000800000000000000000000020000) 
14'h2592 : LOC =         127'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000; // D (0x00001000000000000000000000020000) 
14'h1e81 : LOC =         127'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000; // D (0x00002000000000000000000000020000) 
14'h2bd0 : LOC =         127'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000; // D (0x00004000000000000000000000020000) 
14'h0205 : LOC =         127'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000; // D (0x00008000000000000000000000020000) 
14'h12d8 : LOC =         127'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000; // D (0x00010000000000000000000000020000) 
14'h3362 : LOC =         127'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000; // D (0x00020000000000000000000000020000) 
14'h3361 : LOC =         127'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000; // D (0x00040000000000000000000000020000) 
14'h3367 : LOC =         127'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000; // D (0x00080000000000000000000000020000) 
14'h336b : LOC =         127'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000; // D (0x00100000000000000000000000020000) 
14'h3373 : LOC =         127'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000; // D (0x00200000000000000000000000020000) 
14'h3343 : LOC =         127'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000; // D (0x00400000000000000000000000020000) 
14'h3323 : LOC =         127'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000; // D (0x00800000000000000000000000020000) 
14'h33e3 : LOC =         127'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000; // D (0x01000000000000000000000000020000) 
14'h3263 : LOC =         127'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000; // D (0x02000000000000000000000000020000) 
14'h3163 : LOC =         127'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000; // D (0x04000000000000000000000000020000) 
14'h3763 : LOC =         127'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000; // D (0x08000000000000000000000000020000) 
14'h3b63 : LOC =         127'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000; // D (0x10000000000000000000000000020000) 
14'h2363 : LOC =         127'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000; // D (0x20000000000000000000000000020000) 
14'h1363 : LOC =         127'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000; // D (0x40000000000000000000000000020000) 
14'h25b1 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000; // S (0x00000000000000000000000000040000) 
14'h2da4 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000; // D (0x000000000000000000000000000c0000) 
14'h359b : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000000000000000000; // D (0x00000000000000000000000000140000) 
14'h05e5 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000; // D (0x00000000000000000000000000240000) 
14'h266e : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000000000000000000; // D (0x00000000000000000000000000440000) 
14'h220f : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100001000000000000000000; // D (0x00000000000000000000000000840000) 
14'h2acd : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000001000000000000000000; // D (0x00000000000000000000000001040000) 
14'h3b49 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000001000000000000000000; // D (0x00000000000000000000000002040000) 
14'h1841 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000001000000000000000000; // D (0x00000000000000000000000004040000) 
14'h1d26 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000001000000000000000000; // D (0x00000000000000000000000008040000) 
14'h17e8 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000001000000000000000000; // D (0x00000000000000000000000010040000) 
14'h0274 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000001000000000000000000; // D (0x00000000000000000000000020040000) 
14'h294c : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000001000000000000000000; // D (0x00000000000000000000000040040000) 
14'h3c4b : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000001000000000000000000; // D (0x00000000000000000000000080040000) 
14'h1645 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000001000000000000000000; // D (0x00000000000000000000000100040000) 
14'h012e : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000001000000000000000000; // D (0x00000000000000000000000200040000) 
14'h2ff8 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001000000000000000000; // D (0x00000000000000000000000400040000) 
14'h3123 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000001000000000000000000; // D (0x00000000000000000000000800040000) 
14'h0c95 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000001000000000000000000; // D (0x00000000000000000000001000040000) 
14'h348e : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000001000000000000000000; // D (0x00000000000000000000002000040000) 
14'h07cf : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000001000000000000000000; // D (0x00000000000000000000004000040000) 
14'h223a : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000001000000000000000000; // D (0x00000000000000000000008000040000) 
14'h2aa7 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000001000000000000000000; // D (0x00000000000000000000010000040000) 
14'h3b9d : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000001000000000000000000; // D (0x00000000000000000000020000040000) 
14'h19e9 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000001000000000000000000; // D (0x00000000000000000000040000040000) 
14'h1e76 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000001000000000000000000; // D (0x00000000000000000000080000040000) 
14'h1148 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000001000000000000000000; // D (0x00000000000000000000100000040000) 
14'h0f34 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000001000000000000000000; // D (0x00000000000000000000200000040000) 
14'h33cc : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000001000000000000000000; // D (0x00000000000000000000400000040000) 
14'h094b : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000001000000000000000000; // D (0x00000000000000000000800000040000) 
14'h3f32 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000001000000000000000000; // D (0x00000000000000000001000000040000) 
14'h10b7 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000001000000000000000000; // D (0x00000000000000000002000000040000) 
14'h0cca : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000001000000000000000000; // D (0x00000000000000000004000000040000) 
14'h3430 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000001000000000000000000; // D (0x00000000000000000008000000040000) 
14'h06b3 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000001000000000000000000; // D (0x00000000000000000010000000040000) 
14'h20c2 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000001000000000000000000; // D (0x00000000000000000020000000040000) 
14'h2f57 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000001000000000000000000; // D (0x00000000000000000040000000040000) 
14'h307d : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000001000000000000000000; // D (0x00000000000000000080000000040000) 
14'h0e29 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000000000000; // D (0x00000000000000000100000000040000) 
14'h31f6 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000001000000000000000000; // D (0x00000000000000000200000000040000) 
14'h0d3f : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000001000000000000000000; // D (0x00000000000000000400000000040000) 
14'h37da : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000001000000000000000000; // D (0x00000000000000000800000000040000) 
14'h0167 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000001000000000000000000; // D (0x00000000000000001000000000040000) 
14'h2f6a : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000001000000000000000000; // D (0x00000000000000002000000000040000) 
14'h3007 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000001000000000000000000; // D (0x00000000000000004000000000040000) 
14'h0edd : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000001000000000000000000; // D (0x00000000000000008000000000040000) 
14'h301e : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000001000000000000000000; // D (0x00000000000000010000000000040000) 
14'h0eef : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000001000000000000000000; // D (0x00000000000000020000000000040000) 
14'h307a : LOC =         127'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000001000000000000000000; // D (0x00000000000000040000000000040000) 
14'h0e27 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000001000000000000000000; // D (0x00000000000000080000000000040000) 
14'h31ea : LOC =         127'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000001000000000000000000; // D (0x00000000000000100000000000040000) 
14'h0d07 : LOC =         127'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000001000000000000000000; // D (0x00000000000000200000000000040000) 
14'h37aa : LOC =         127'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000001000000000000000000; // D (0x00000000000000400000000000040000) 
14'h0187 : LOC =         127'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000001000000000000000000; // D (0x00000000000000800000000000040000) 
14'h2eaa : LOC =         127'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000001000000000000000000; // D (0x00000000000001000000000000040000) 
14'h3387 : LOC =         127'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000001000000000000000000; // D (0x00000000000002000000000000040000) 
14'h09dd : LOC =         127'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000001000000000000000000; // D (0x00000000000004000000000000040000) 
14'h3e1e : LOC =         127'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000001000000000000000000; // D (0x00000000000008000000000000040000) 
14'h12ef : LOC =         127'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000001000000000000000000; // D (0x00000000000010000000000000040000) 
14'h087a : LOC =         127'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000001000000000000000000; // D (0x00000000000020000000000000040000) 
14'h3d50 : LOC =         127'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000001000000000000000000; // D (0x00000000000040000000000000040000) 
14'h1473 : LOC =         127'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000001000000000000000000; // D (0x00000000000080000000000000040000) 
14'h0542 : LOC =         127'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000001000000000000000000; // D (0x00000000000100000000000000040000) 
14'h2720 : LOC =         127'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000001000000000000000000; // D (0x00000000000200000000000000040000) 
14'h2093 : LOC =         127'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000001000000000000000000; // D (0x00000000000400000000000000040000) 
14'h2ff5 : LOC =         127'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000001000000000000000000; // D (0x00000000000800000000000000040000) 
14'h3139 : LOC =         127'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000001000000000000000000; // D (0x00000000001000000000000000040000) 
14'h0ca1 : LOC =         127'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000001000000000000000000; // D (0x00000000002000000000000000040000) 
14'h34e6 : LOC =         127'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000001000000000000000000; // D (0x00000000004000000000000000040000) 
14'h071f : LOC =         127'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000001000000000000000000; // D (0x00000000008000000000000000040000) 
14'h239a : LOC =         127'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000001000000000000000000; // D (0x00000000010000000000000000040000) 
14'h29e7 : LOC =         127'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000001000000000000000000; // D (0x00000000020000000000000000040000) 
14'h3d1d : LOC =         127'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000; // D (0x00000000040000000000000000040000) 
14'h14e9 : LOC =         127'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000; // D (0x00000000080000000000000000040000) 
14'h0476 : LOC =         127'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000; // D (0x00000000100000000000000000040000) 
14'h2548 : LOC =         127'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000; // D (0x00000000200000000000000000040000) 
14'h2443 : LOC =         127'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000; // D (0x00000000400000000000000000040000) 
14'h2655 : LOC =         127'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000; // D (0x00000000800000000000000000040000) 
14'h2279 : LOC =         127'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000; // D (0x00000001000000000000000000040000) 
14'h2a21 : LOC =         127'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000; // D (0x00000002000000000000000000040000) 
14'h3a91 : LOC =         127'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000; // D (0x00000004000000000000000000040000) 
14'h1bf1 : LOC =         127'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000; // D (0x00000008000000000000000000040000) 
14'h1a46 : LOC =         127'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000; // D (0x00000010000000000000000000040000) 
14'h1928 : LOC =         127'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000; // D (0x00000020000000000000000000040000) 
14'h1ff4 : LOC =         127'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000; // D (0x00000040000000000000000000040000) 
14'h124c : LOC =         127'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000; // D (0x00000080000000000000000000040000) 
14'h093c : LOC =         127'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000; // D (0x00000100000000000000000000040000) 
14'h3fdc : LOC =         127'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000; // D (0x00000200000000000000000000040000) 
14'h116b : LOC =         127'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000; // D (0x00000400000000000000000000040000) 
14'h0f72 : LOC =         127'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000; // D (0x00000800000000000000000000040000) 
14'h3340 : LOC =         127'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000; // D (0x00001000000000000000000000040000) 
14'h0853 : LOC =         127'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000; // D (0x00002000000000000000000000040000) 
14'h3d02 : LOC =         127'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000; // D (0x00004000000000000000000000040000) 
14'h14d7 : LOC =         127'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000; // D (0x00008000000000000000000000040000) 
14'h040a : LOC =         127'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000; // D (0x00010000000000000000000000040000) 
14'h25b0 : LOC =         127'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000; // D (0x00020000000000000000000000040000) 
14'h25b3 : LOC =         127'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000; // D (0x00040000000000000000000000040000) 
14'h25b5 : LOC =         127'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000; // D (0x00080000000000000000000000040000) 
14'h25b9 : LOC =         127'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000; // D (0x00100000000000000000000000040000) 
14'h25a1 : LOC =         127'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000; // D (0x00200000000000000000000000040000) 
14'h2591 : LOC =         127'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000; // D (0x00400000000000000000000000040000) 
14'h25f1 : LOC =         127'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000; // D (0x00800000000000000000000000040000) 
14'h2531 : LOC =         127'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000; // D (0x01000000000000000000000000040000) 
14'h24b1 : LOC =         127'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000; // D (0x02000000000000000000000000040000) 
14'h27b1 : LOC =         127'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000; // D (0x04000000000000000000000000040000) 
14'h21b1 : LOC =         127'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000; // D (0x08000000000000000000000000040000) 
14'h2db1 : LOC =         127'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000; // D (0x10000000000000000000000000040000) 
14'h35b1 : LOC =         127'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000; // D (0x20000000000000000000000000040000) 
14'h05b1 : LOC =         127'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000; // D (0x40000000000000000000000000040000) 
14'h0815 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000; // S (0x00000000000000000000000000080000) 
14'h183f : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000; // D (0x00000000000000000000000000180000) 
14'h2841 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000000000000000000; // D (0x00000000000000000000000000280000) 
14'h0bca : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000; // D (0x00000000000000000000000000480000) 
14'h0fab : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010000000000000000000; // D (0x00000000000000000000000000880000) 
14'h0769 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000010000000000000000000; // D (0x00000000000000000000000001080000) 
14'h16ed : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000010000000000000000000; // D (0x00000000000000000000000002080000) 
14'h35e5 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000010000000000000000000; // D (0x00000000000000000000000004080000) 
14'h3082 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000010000000000000000000; // D (0x00000000000000000000000008080000) 
14'h3a4c : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000010000000000000000000; // D (0x00000000000000000000000010080000) 
14'h2fd0 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000010000000000000000000; // D (0x00000000000000000000000020080000) 
14'h04e8 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000010000000000000000000; // D (0x00000000000000000000000040080000) 
14'h11ef : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000010000000000000000000; // D (0x00000000000000000000000080080000) 
14'h3be1 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000010000000000000000000; // D (0x00000000000000000000000100080000) 
14'h2c8a : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000010000000000000000000; // D (0x00000000000000000000000200080000) 
14'h025c : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000010000000000000000000; // D (0x00000000000000000000000400080000) 
14'h1c87 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000010000000000000000000; // D (0x00000000000000000000000800080000) 
14'h2131 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000010000000000000000000; // D (0x00000000000000000000001000080000) 
14'h192a : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000010000000000000000000; // D (0x00000000000000000000002000080000) 
14'h2a6b : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000010000000000000000000; // D (0x00000000000000000000004000080000) 
14'h0f9e : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000010000000000000000000; // D (0x00000000000000000000008000080000) 
14'h0703 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000010000000000000000000; // D (0x00000000000000000000010000080000) 
14'h1639 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000010000000000000000000; // D (0x00000000000000000000020000080000) 
14'h344d : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000010000000000000000000; // D (0x00000000000000000000040000080000) 
14'h33d2 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000010000000000000000000; // D (0x00000000000000000000080000080000) 
14'h3cec : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000010000000000000000000; // D (0x00000000000000000000100000080000) 
14'h2290 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000010000000000000000000; // D (0x00000000000000000000200000080000) 
14'h1e68 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000010000000000000000000; // D (0x00000000000000000000400000080000) 
14'h24ef : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000010000000000000000000; // D (0x00000000000000000000800000080000) 
14'h1296 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000010000000000000000000; // D (0x00000000000000000001000000080000) 
14'h3d13 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000010000000000000000000; // D (0x00000000000000000002000000080000) 
14'h216e : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000010000000000000000000; // D (0x00000000000000000004000000080000) 
14'h1994 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000010000000000000000000; // D (0x00000000000000000008000000080000) 
14'h2b17 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000010000000000000000000; // D (0x00000000000000000010000000080000) 
14'h0d66 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000010000000000000000000; // D (0x00000000000000000020000000080000) 
14'h02f3 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000010000000000000000000; // D (0x00000000000000000040000000080000) 
14'h1dd9 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000010000000000000000000; // D (0x00000000000000000080000000080000) 
14'h238d : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000010000000000000000000; // D (0x00000000000000000100000000080000) 
14'h1c52 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000010000000000000000000; // D (0x00000000000000000200000000080000) 
14'h209b : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000010000000000000000000; // D (0x00000000000000000400000000080000) 
14'h1a7e : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000010000000000000000000; // D (0x00000000000000000800000000080000) 
14'h2cc3 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000010000000000000000000; // D (0x00000000000000001000000000080000) 
14'h02ce : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000010000000000000000000; // D (0x00000000000000002000000000080000) 
14'h1da3 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000010000000000000000000; // D (0x00000000000000004000000000080000) 
14'h2379 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000010000000000000000000; // D (0x00000000000000008000000000080000) 
14'h1dba : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000010000000000000000000; // D (0x00000000000000010000000000080000) 
14'h234b : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000010000000000000000000; // D (0x00000000000000020000000000080000) 
14'h1dde : LOC =         127'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000010000000000000000000; // D (0x00000000000000040000000000080000) 
14'h2383 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000010000000000000000000; // D (0x00000000000000080000000000080000) 
14'h1c4e : LOC =         127'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000010000000000000000000; // D (0x00000000000000100000000000080000) 
14'h20a3 : LOC =         127'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000010000000000000000000; // D (0x00000000000000200000000000080000) 
14'h1a0e : LOC =         127'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000010000000000000000000; // D (0x00000000000000400000000000080000) 
14'h2c23 : LOC =         127'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000010000000000000000000; // D (0x00000000000000800000000000080000) 
14'h030e : LOC =         127'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000010000000000000000000; // D (0x00000000000001000000000000080000) 
14'h1e23 : LOC =         127'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000010000000000000000000; // D (0x00000000000002000000000000080000) 
14'h2479 : LOC =         127'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000010000000000000000000; // D (0x00000000000004000000000000080000) 
14'h13ba : LOC =         127'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000010000000000000000000; // D (0x00000000000008000000000000080000) 
14'h3f4b : LOC =         127'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000010000000000000000000; // D (0x00000000000010000000000000080000) 
14'h25de : LOC =         127'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000010000000000000000000; // D (0x00000000000020000000000000080000) 
14'h10f4 : LOC =         127'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000010000000000000000000; // D (0x00000000000040000000000000080000) 
14'h39d7 : LOC =         127'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000010000000000000000000; // D (0x00000000000080000000000000080000) 
14'h28e6 : LOC =         127'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000010000000000000000000; // D (0x00000000000100000000000000080000) 
14'h0a84 : LOC =         127'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000010000000000000000000; // D (0x00000000000200000000000000080000) 
14'h0d37 : LOC =         127'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000010000000000000000000; // D (0x00000000000400000000000000080000) 
14'h0251 : LOC =         127'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000010000000000000000000; // D (0x00000000000800000000000000080000) 
14'h1c9d : LOC =         127'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000010000000000000000000; // D (0x00000000001000000000000000080000) 
14'h2105 : LOC =         127'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000010000000000000000000; // D (0x00000000002000000000000000080000) 
14'h1942 : LOC =         127'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000010000000000000000000; // D (0x00000000004000000000000000080000) 
14'h2abb : LOC =         127'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000010000000000000000000; // D (0x00000000008000000000000000080000) 
14'h0e3e : LOC =         127'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000010000000000000000000; // D (0x00000000010000000000000000080000) 
14'h0443 : LOC =         127'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000010000000000000000000; // D (0x00000000020000000000000000080000) 
14'h10b9 : LOC =         127'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000; // D (0x00000000040000000000000000080000) 
14'h394d : LOC =         127'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000; // D (0x00000000080000000000000000080000) 
14'h29d2 : LOC =         127'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000; // D (0x00000000100000000000000000080000) 
14'h08ec : LOC =         127'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000; // D (0x00000000200000000000000000080000) 
14'h09e7 : LOC =         127'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000; // D (0x00000000400000000000000000080000) 
14'h0bf1 : LOC =         127'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000; // D (0x00000000800000000000000000080000) 
14'h0fdd : LOC =         127'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000; // D (0x00000001000000000000000000080000) 
14'h0785 : LOC =         127'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000; // D (0x00000002000000000000000000080000) 
14'h1735 : LOC =         127'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000; // D (0x00000004000000000000000000080000) 
14'h3655 : LOC =         127'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000; // D (0x00000008000000000000000000080000) 
14'h37e2 : LOC =         127'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000; // D (0x00000010000000000000000000080000) 
14'h348c : LOC =         127'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000; // D (0x00000020000000000000000000080000) 
14'h3250 : LOC =         127'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000; // D (0x00000040000000000000000000080000) 
14'h3fe8 : LOC =         127'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000; // D (0x00000080000000000000000000080000) 
14'h2498 : LOC =         127'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000; // D (0x00000100000000000000000000080000) 
14'h1278 : LOC =         127'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000; // D (0x00000200000000000000000000080000) 
14'h3ccf : LOC =         127'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000; // D (0x00000400000000000000000000080000) 
14'h22d6 : LOC =         127'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000; // D (0x00000800000000000000000000080000) 
14'h1ee4 : LOC =         127'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000; // D (0x00001000000000000000000000080000) 
14'h25f7 : LOC =         127'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000; // D (0x00002000000000000000000000080000) 
14'h10a6 : LOC =         127'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000; // D (0x00004000000000000000000000080000) 
14'h3973 : LOC =         127'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000; // D (0x00008000000000000000000000080000) 
14'h29ae : LOC =         127'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000; // D (0x00010000000000000000000000080000) 
14'h0814 : LOC =         127'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000; // D (0x00020000000000000000000000080000) 
14'h0817 : LOC =         127'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000; // D (0x00040000000000000000000000080000) 
14'h0811 : LOC =         127'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000; // D (0x00080000000000000000000000080000) 
14'h081d : LOC =         127'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000; // D (0x00100000000000000000000000080000) 
14'h0805 : LOC =         127'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000; // D (0x00200000000000000000000000080000) 
14'h0835 : LOC =         127'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000; // D (0x00400000000000000000000000080000) 
14'h0855 : LOC =         127'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000; // D (0x00800000000000000000000000080000) 
14'h0895 : LOC =         127'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000; // D (0x01000000000000000000000000080000) 
14'h0915 : LOC =         127'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000; // D (0x02000000000000000000000000080000) 
14'h0a15 : LOC =         127'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000; // D (0x04000000000000000000000000080000) 
14'h0c15 : LOC =         127'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000; // D (0x08000000000000000000000000080000) 
14'h0015 : LOC =         127'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000; // D (0x10000000000000000000000000080000) 
14'h1815 : LOC =         127'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000; // D (0x20000000000000000000000000080000) 
14'h2815 : LOC =         127'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000; // D (0x40000000000000000000000000080000) 
14'h102a : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000; // S (0x00000000000000000000000000100000) 
14'h307e : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000; // D (0x00000000000000000000000000300000) 
14'h13f5 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000; // D (0x00000000000000000000000000500000) 
14'h1794 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000; // D (0x00000000000000000000000000900000) 
14'h1f56 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000100000000000000000000; // D (0x00000000000000000000000001100000) 
14'h0ed2 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000100000000000000000000; // D (0x00000000000000000000000002100000) 
14'h2dda : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000100000000000000000000; // D (0x00000000000000000000000004100000) 
14'h28bd : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000100000000000000000000; // D (0x00000000000000000000000008100000) 
14'h2273 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000100000000000000000000; // D (0x00000000000000000000000010100000) 
14'h37ef : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000100000000000000000000; // D (0x00000000000000000000000020100000) 
14'h1cd7 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000100000000000000000000; // D (0x00000000000000000000000040100000) 
14'h09d0 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000100000000000000000000; // D (0x00000000000000000000000080100000) 
14'h23de : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000100000000000000000000; // D (0x00000000000000000000000100100000) 
14'h34b5 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000100000000000000000000; // D (0x00000000000000000000000200100000) 
14'h1a63 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000100000000000000000000; // D (0x00000000000000000000000400100000) 
14'h04b8 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000100000000000000000000; // D (0x00000000000000000000000800100000) 
14'h390e : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000100000000000000000000; // D (0x00000000000000000000001000100000) 
14'h0115 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000100000000000000000000; // D (0x00000000000000000000002000100000) 
14'h3254 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000100000000000000000000; // D (0x00000000000000000000004000100000) 
14'h17a1 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000100000000000000000000; // D (0x00000000000000000000008000100000) 
14'h1f3c : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000100000000000000000000; // D (0x00000000000000000000010000100000) 
14'h0e06 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000100000000000000000000; // D (0x00000000000000000000020000100000) 
14'h2c72 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000100000000000000000000; // D (0x00000000000000000000040000100000) 
14'h2bed : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000100000000000000000000; // D (0x00000000000000000000080000100000) 
14'h24d3 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000100000000000000000000; // D (0x00000000000000000000100000100000) 
14'h3aaf : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000100000000000000000000; // D (0x00000000000000000000200000100000) 
14'h0657 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000100000000000000000000; // D (0x00000000000000000000400000100000) 
14'h3cd0 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000100000000000000000000; // D (0x00000000000000000000800000100000) 
14'h0aa9 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000100000000000000000000; // D (0x00000000000000000001000000100000) 
14'h252c : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000100000000000000000000; // D (0x00000000000000000002000000100000) 
14'h3951 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000100000000000000000000; // D (0x00000000000000000004000000100000) 
14'h01ab : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000100000000000000000000; // D (0x00000000000000000008000000100000) 
14'h3328 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000100000000000000000000; // D (0x00000000000000000010000000100000) 
14'h1559 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000100000000000000000000; // D (0x00000000000000000020000000100000) 
14'h1acc : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000100000000000000000000; // D (0x00000000000000000040000000100000) 
14'h05e6 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000100000000000000000000; // D (0x00000000000000000080000000100000) 
14'h3bb2 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000100000000000000000000; // D (0x00000000000000000100000000100000) 
14'h046d : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000100000000000000000000; // D (0x00000000000000000200000000100000) 
14'h38a4 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000100000000000000000000; // D (0x00000000000000000400000000100000) 
14'h0241 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000100000000000000000000; // D (0x00000000000000000800000000100000) 
14'h34fc : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000100000000000000000000; // D (0x00000000000000001000000000100000) 
14'h1af1 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000100000000000000000000; // D (0x00000000000000002000000000100000) 
14'h059c : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000100000000000000000000; // D (0x00000000000000004000000000100000) 
14'h3b46 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000100000000000000000000; // D (0x00000000000000008000000000100000) 
14'h0585 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000100000000000000000000; // D (0x00000000000000010000000000100000) 
14'h3b74 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000100000000000000000000; // D (0x00000000000000020000000000100000) 
14'h05e1 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000100000000000000000000; // D (0x00000000000000040000000000100000) 
14'h3bbc : LOC =         127'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000100000000000000000000; // D (0x00000000000000080000000000100000) 
14'h0471 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000100000000000000000000; // D (0x00000000000000100000000000100000) 
14'h389c : LOC =         127'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000100000000000000000000; // D (0x00000000000000200000000000100000) 
14'h0231 : LOC =         127'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000100000000000000000000; // D (0x00000000000000400000000000100000) 
14'h341c : LOC =         127'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000100000000000000000000; // D (0x00000000000000800000000000100000) 
14'h1b31 : LOC =         127'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000100000000000000000000; // D (0x00000000000001000000000000100000) 
14'h061c : LOC =         127'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000100000000000000000000; // D (0x00000000000002000000000000100000) 
14'h3c46 : LOC =         127'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000100000000000000000000; // D (0x00000000000004000000000000100000) 
14'h0b85 : LOC =         127'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000100000000000000000000; // D (0x00000000000008000000000000100000) 
14'h2774 : LOC =         127'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000100000000000000000000; // D (0x00000000000010000000000000100000) 
14'h3de1 : LOC =         127'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000100000000000000000000; // D (0x00000000000020000000000000100000) 
14'h08cb : LOC =         127'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000100000000000000000000; // D (0x00000000000040000000000000100000) 
14'h21e8 : LOC =         127'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000100000000000000000000; // D (0x00000000000080000000000000100000) 
14'h30d9 : LOC =         127'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000100000000000000000000; // D (0x00000000000100000000000000100000) 
14'h12bb : LOC =         127'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000100000000000000000000; // D (0x00000000000200000000000000100000) 
14'h1508 : LOC =         127'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000100000000000000000000; // D (0x00000000000400000000000000100000) 
14'h1a6e : LOC =         127'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000100000000000000000000; // D (0x00000000000800000000000000100000) 
14'h04a2 : LOC =         127'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000100000000000000000000; // D (0x00000000001000000000000000100000) 
14'h393a : LOC =         127'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000100000000000000000000; // D (0x00000000002000000000000000100000) 
14'h017d : LOC =         127'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000100000000000000000000; // D (0x00000000004000000000000000100000) 
14'h3284 : LOC =         127'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000100000000000000000000; // D (0x00000000008000000000000000100000) 
14'h1601 : LOC =         127'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000100000000000000000000; // D (0x00000000010000000000000000100000) 
14'h1c7c : LOC =         127'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000100000000000000000000; // D (0x00000000020000000000000000100000) 
14'h0886 : LOC =         127'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000; // D (0x00000000040000000000000000100000) 
14'h2172 : LOC =         127'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000; // D (0x00000000080000000000000000100000) 
14'h31ed : LOC =         127'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000; // D (0x00000000100000000000000000100000) 
14'h10d3 : LOC =         127'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000; // D (0x00000000200000000000000000100000) 
14'h11d8 : LOC =         127'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000; // D (0x00000000400000000000000000100000) 
14'h13ce : LOC =         127'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000; // D (0x00000000800000000000000000100000) 
14'h17e2 : LOC =         127'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000; // D (0x00000001000000000000000000100000) 
14'h1fba : LOC =         127'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000; // D (0x00000002000000000000000000100000) 
14'h0f0a : LOC =         127'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000; // D (0x00000004000000000000000000100000) 
14'h2e6a : LOC =         127'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000; // D (0x00000008000000000000000000100000) 
14'h2fdd : LOC =         127'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000; // D (0x00000010000000000000000000100000) 
14'h2cb3 : LOC =         127'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000; // D (0x00000020000000000000000000100000) 
14'h2a6f : LOC =         127'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000; // D (0x00000040000000000000000000100000) 
14'h27d7 : LOC =         127'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000; // D (0x00000080000000000000000000100000) 
14'h3ca7 : LOC =         127'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000; // D (0x00000100000000000000000000100000) 
14'h0a47 : LOC =         127'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000; // D (0x00000200000000000000000000100000) 
14'h24f0 : LOC =         127'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000; // D (0x00000400000000000000000000100000) 
14'h3ae9 : LOC =         127'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000; // D (0x00000800000000000000000000100000) 
14'h06db : LOC =         127'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000; // D (0x00001000000000000000000000100000) 
14'h3dc8 : LOC =         127'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000; // D (0x00002000000000000000000000100000) 
14'h0899 : LOC =         127'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000; // D (0x00004000000000000000000000100000) 
14'h214c : LOC =         127'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000; // D (0x00008000000000000000000000100000) 
14'h3191 : LOC =         127'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000; // D (0x00010000000000000000000000100000) 
14'h102b : LOC =         127'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000; // D (0x00020000000000000000000000100000) 
14'h1028 : LOC =         127'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000; // D (0x00040000000000000000000000100000) 
14'h102e : LOC =         127'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000; // D (0x00080000000000000000000000100000) 
14'h1022 : LOC =         127'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000; // D (0x00100000000000000000000000100000) 
14'h103a : LOC =         127'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000; // D (0x00200000000000000000000000100000) 
14'h100a : LOC =         127'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000; // D (0x00400000000000000000000000100000) 
14'h106a : LOC =         127'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000; // D (0x00800000000000000000000000100000) 
14'h10aa : LOC =         127'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000; // D (0x01000000000000000000000000100000) 
14'h112a : LOC =         127'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000; // D (0x02000000000000000000000000100000) 
14'h122a : LOC =         127'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000; // D (0x04000000000000000000000000100000) 
14'h142a : LOC =         127'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000; // D (0x08000000000000000000000000100000) 
14'h182a : LOC =         127'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000; // D (0x10000000000000000000000000100000) 
14'h002a : LOC =         127'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000; // D (0x20000000000000000000000000100000) 
14'h302a : LOC =         127'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000; // D (0x40000000000000000000000000100000) 
14'h2054 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000; // S (0x00000000000000000000000000200000) 
14'h238b : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000; // D (0x00000000000000000000000000600000) 
14'h27ea : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000000000000000000000; // D (0x00000000000000000000000000a00000) 
14'h2f28 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000000; // D (0x00000000000000000000000001200000) 
14'h3eac : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000000000000000000000; // D (0x00000000000000000000000002200000) 
14'h1da4 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100001000000000000000000000; // D (0x00000000000000000000000004200000) 
14'h18c3 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000001000000000000000000000; // D (0x00000000000000000000000008200000) 
14'h120d : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000001000000000000000000000; // D (0x00000000000000000000000010200000) 
14'h0791 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000001000000000000000000000; // D (0x00000000000000000000000020200000) 
14'h2ca9 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000001000000000000000000000; // D (0x00000000000000000000000040200000) 
14'h39ae : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000001000000000000000000000; // D (0x00000000000000000000000080200000) 
14'h13a0 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000001000000000000000000000; // D (0x00000000000000000000000100200000) 
14'h04cb : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000001000000000000000000000; // D (0x00000000000000000000000200200000) 
14'h2a1d : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000001000000000000000000000; // D (0x00000000000000000000000400200000) 
14'h34c6 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000001000000000000000000000; // D (0x00000000000000000000000800200000) 
14'h0970 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000001000000000000000000000; // D (0x00000000000000000000001000200000) 
14'h316b : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001000000000000000000000; // D (0x00000000000000000000002000200000) 
14'h022a : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000001000000000000000000000; // D (0x00000000000000000000004000200000) 
14'h27df : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000001000000000000000000000; // D (0x00000000000000000000008000200000) 
14'h2f42 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000001000000000000000000000; // D (0x00000000000000000000010000200000) 
14'h3e78 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000001000000000000000000000; // D (0x00000000000000000000020000200000) 
14'h1c0c : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000001000000000000000000000; // D (0x00000000000000000000040000200000) 
14'h1b93 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000001000000000000000000000; // D (0x00000000000000000000080000200000) 
14'h14ad : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000001000000000000000000000; // D (0x00000000000000000000100000200000) 
14'h0ad1 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000001000000000000000000000; // D (0x00000000000000000000200000200000) 
14'h3629 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000001000000000000000000000; // D (0x00000000000000000000400000200000) 
14'h0cae : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000001000000000000000000000; // D (0x00000000000000000000800000200000) 
14'h3ad7 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000001000000000000000000000; // D (0x00000000000000000001000000200000) 
14'h1552 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000001000000000000000000000; // D (0x00000000000000000002000000200000) 
14'h092f : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000001000000000000000000000; // D (0x00000000000000000004000000200000) 
14'h31d5 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000001000000000000000000000; // D (0x00000000000000000008000000200000) 
14'h0356 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000001000000000000000000000; // D (0x00000000000000000010000000200000) 
14'h2527 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000001000000000000000000000; // D (0x00000000000000000020000000200000) 
14'h2ab2 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000001000000000000000000000; // D (0x00000000000000000040000000200000) 
14'h3598 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000001000000000000000000000; // D (0x00000000000000000080000000200000) 
14'h0bcc : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000001000000000000000000000; // D (0x00000000000000000100000000200000) 
14'h3413 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000001000000000000000000000; // D (0x00000000000000000200000000200000) 
14'h08da : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000001000000000000000000000; // D (0x00000000000000000400000000200000) 
14'h323f : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000000000000000; // D (0x00000000000000000800000000200000) 
14'h0482 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000001000000000000000000000; // D (0x00000000000000001000000000200000) 
14'h2a8f : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000001000000000000000000000; // D (0x00000000000000002000000000200000) 
14'h35e2 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000001000000000000000000000; // D (0x00000000000000004000000000200000) 
14'h0b38 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000001000000000000000000000; // D (0x00000000000000008000000000200000) 
14'h35fb : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000001000000000000000000000; // D (0x00000000000000010000000000200000) 
14'h0b0a : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000001000000000000000000000; // D (0x00000000000000020000000000200000) 
14'h359f : LOC =         127'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000001000000000000000000000; // D (0x00000000000000040000000000200000) 
14'h0bc2 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000001000000000000000000000; // D (0x00000000000000080000000000200000) 
14'h340f : LOC =         127'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000001000000000000000000000; // D (0x00000000000000100000000000200000) 
14'h08e2 : LOC =         127'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000001000000000000000000000; // D (0x00000000000000200000000000200000) 
14'h324f : LOC =         127'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000001000000000000000000000; // D (0x00000000000000400000000000200000) 
14'h0462 : LOC =         127'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000001000000000000000000000; // D (0x00000000000000800000000000200000) 
14'h2b4f : LOC =         127'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000001000000000000000000000; // D (0x00000000000001000000000000200000) 
14'h3662 : LOC =         127'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000001000000000000000000000; // D (0x00000000000002000000000000200000) 
14'h0c38 : LOC =         127'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000001000000000000000000000; // D (0x00000000000004000000000000200000) 
14'h3bfb : LOC =         127'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000001000000000000000000000; // D (0x00000000000008000000000000200000) 
14'h170a : LOC =         127'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000001000000000000000000000; // D (0x00000000000010000000000000200000) 
14'h0d9f : LOC =         127'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000001000000000000000000000; // D (0x00000000000020000000000000200000) 
14'h38b5 : LOC =         127'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000001000000000000000000000; // D (0x00000000000040000000000000200000) 
14'h1196 : LOC =         127'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000001000000000000000000000; // D (0x00000000000080000000000000200000) 
14'h00a7 : LOC =         127'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000001000000000000000000000; // D (0x00000000000100000000000000200000) 
14'h22c5 : LOC =         127'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000001000000000000000000000; // D (0x00000000000200000000000000200000) 
14'h2576 : LOC =         127'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000001000000000000000000000; // D (0x00000000000400000000000000200000) 
14'h2a10 : LOC =         127'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000001000000000000000000000; // D (0x00000000000800000000000000200000) 
14'h34dc : LOC =         127'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000001000000000000000000000; // D (0x00000000001000000000000000200000) 
14'h0944 : LOC =         127'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000001000000000000000000000; // D (0x00000000002000000000000000200000) 
14'h3103 : LOC =         127'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000001000000000000000000000; // D (0x00000000004000000000000000200000) 
14'h02fa : LOC =         127'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000001000000000000000000000; // D (0x00000000008000000000000000200000) 
14'h267f : LOC =         127'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000001000000000000000000000; // D (0x00000000010000000000000000200000) 
14'h2c02 : LOC =         127'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000001000000000000000000000; // D (0x00000000020000000000000000200000) 
14'h38f8 : LOC =         127'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000; // D (0x00000000040000000000000000200000) 
14'h110c : LOC =         127'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000; // D (0x00000000080000000000000000200000) 
14'h0193 : LOC =         127'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000; // D (0x00000000100000000000000000200000) 
14'h20ad : LOC =         127'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000; // D (0x00000000200000000000000000200000) 
14'h21a6 : LOC =         127'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000; // D (0x00000000400000000000000000200000) 
14'h23b0 : LOC =         127'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000; // D (0x00000000800000000000000000200000) 
14'h279c : LOC =         127'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000; // D (0x00000001000000000000000000200000) 
14'h2fc4 : LOC =         127'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000; // D (0x00000002000000000000000000200000) 
14'h3f74 : LOC =         127'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000; // D (0x00000004000000000000000000200000) 
14'h1e14 : LOC =         127'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000; // D (0x00000008000000000000000000200000) 
14'h1fa3 : LOC =         127'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000; // D (0x00000010000000000000000000200000) 
14'h1ccd : LOC =         127'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000; // D (0x00000020000000000000000000200000) 
14'h1a11 : LOC =         127'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000; // D (0x00000040000000000000000000200000) 
14'h17a9 : LOC =         127'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000; // D (0x00000080000000000000000000200000) 
14'h0cd9 : LOC =         127'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000; // D (0x00000100000000000000000000200000) 
14'h3a39 : LOC =         127'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000; // D (0x00000200000000000000000000200000) 
14'h148e : LOC =         127'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000; // D (0x00000400000000000000000000200000) 
14'h0a97 : LOC =         127'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000; // D (0x00000800000000000000000000200000) 
14'h36a5 : LOC =         127'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000; // D (0x00001000000000000000000000200000) 
14'h0db6 : LOC =         127'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000; // D (0x00002000000000000000000000200000) 
14'h38e7 : LOC =         127'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000; // D (0x00004000000000000000000000200000) 
14'h1132 : LOC =         127'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000; // D (0x00008000000000000000000000200000) 
14'h01ef : LOC =         127'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000; // D (0x00010000000000000000000000200000) 
14'h2055 : LOC =         127'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000; // D (0x00020000000000000000000000200000) 
14'h2056 : LOC =         127'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000; // D (0x00040000000000000000000000200000) 
14'h2050 : LOC =         127'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000; // D (0x00080000000000000000000000200000) 
14'h205c : LOC =         127'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000; // D (0x00100000000000000000000000200000) 
14'h2044 : LOC =         127'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000; // D (0x00200000000000000000000000200000) 
14'h2074 : LOC =         127'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000; // D (0x00400000000000000000000000200000) 
14'h2014 : LOC =         127'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000; // D (0x00800000000000000000000000200000) 
14'h20d4 : LOC =         127'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000; // D (0x01000000000000000000000000200000) 
14'h2154 : LOC =         127'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000; // D (0x02000000000000000000000000200000) 
14'h2254 : LOC =         127'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000; // D (0x04000000000000000000000000200000) 
14'h2454 : LOC =         127'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000; // D (0x08000000000000000000000000200000) 
14'h2854 : LOC =         127'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000; // D (0x10000000000000000000000000200000) 
14'h3054 : LOC =         127'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000; // D (0x20000000000000000000000000200000) 
14'h0054 : LOC =         127'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000; // D (0x40000000000000000000000000200000) 
14'h03df : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000; // S (0x00000000000000000000000000400000) 
14'h0461 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000; // D (0x00000000000000000000000000c00000) 
14'h0ca3 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000000000000000000000; // D (0x00000000000000000000000001400000) 
14'h1d27 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000; // D (0x00000000000000000000000002400000) 
14'h3e2f : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010000000000000000000000; // D (0x00000000000000000000000004400000) 
14'h3b48 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000010000000000000000000000; // D (0x00000000000000000000000008400000) 
14'h3186 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000010000000000000000000000; // D (0x00000000000000000000000010400000) 
14'h241a : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000010000000000000000000000; // D (0x00000000000000000000000020400000) 
14'h0f22 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000010000000000000000000000; // D (0x00000000000000000000000040400000) 
14'h1a25 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000010000000000000000000000; // D (0x00000000000000000000000080400000) 
14'h302b : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000010000000000000000000000; // D (0x00000000000000000000000100400000) 
14'h2740 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000010000000000000000000000; // D (0x00000000000000000000000200400000) 
14'h0996 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000010000000000000000000000; // D (0x00000000000000000000000400400000) 
14'h174d : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000010000000000000000000000; // D (0x00000000000000000000000800400000) 
14'h2afb : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000010000000000000000000000; // D (0x00000000000000000000001000400000) 
14'h12e0 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000010000000000000000000000; // D (0x00000000000000000000002000400000) 
14'h21a1 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000010000000000000000000000; // D (0x00000000000000000000004000400000) 
14'h0454 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000010000000000000000000000; // D (0x00000000000000000000008000400000) 
14'h0cc9 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000010000000000000000000000; // D (0x00000000000000000000010000400000) 
14'h1df3 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000010000000000000000000000; // D (0x00000000000000000000020000400000) 
14'h3f87 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000010000000000000000000000; // D (0x00000000000000000000040000400000) 
14'h3818 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000010000000000000000000000; // D (0x00000000000000000000080000400000) 
14'h3726 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000010000000000000000000000; // D (0x00000000000000000000100000400000) 
14'h295a : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000010000000000000000000000; // D (0x00000000000000000000200000400000) 
14'h15a2 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000010000000000000000000000; // D (0x00000000000000000000400000400000) 
14'h2f25 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000010000000000000000000000; // D (0x00000000000000000000800000400000) 
14'h195c : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000010000000000000000000000; // D (0x00000000000000000001000000400000) 
14'h36d9 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000010000000000000000000000; // D (0x00000000000000000002000000400000) 
14'h2aa4 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000010000000000000000000000; // D (0x00000000000000000004000000400000) 
14'h125e : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000010000000000000000000000; // D (0x00000000000000000008000000400000) 
14'h20dd : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000010000000000000000000000; // D (0x00000000000000000010000000400000) 
14'h06ac : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000010000000000000000000000; // D (0x00000000000000000020000000400000) 
14'h0939 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000010000000000000000000000; // D (0x00000000000000000040000000400000) 
14'h1613 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000010000000000000000000000; // D (0x00000000000000000080000000400000) 
14'h2847 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000; // D (0x00000000000000000100000000400000) 
14'h1798 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000010000000000000000000000; // D (0x00000000000000000200000000400000) 
14'h2b51 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000010000000000000000000000; // D (0x00000000000000000400000000400000) 
14'h11b4 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000010000000000000000000000; // D (0x00000000000000000800000000400000) 
14'h2709 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000010000000000000000000000; // D (0x00000000000000001000000000400000) 
14'h0904 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000010000000000000000000000; // D (0x00000000000000002000000000400000) 
14'h1669 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000010000000000000000000000; // D (0x00000000000000004000000000400000) 
14'h28b3 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000010000000000000000000000; // D (0x00000000000000008000000000400000) 
14'h1670 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000010000000000000000000000; // D (0x00000000000000010000000000400000) 
14'h2881 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000010000000000000000000000; // D (0x00000000000000020000000000400000) 
14'h1614 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000010000000000000000000000; // D (0x00000000000000040000000000400000) 
14'h2849 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000010000000000000000000000; // D (0x00000000000000080000000000400000) 
14'h1784 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000010000000000000000000000; // D (0x00000000000000100000000000400000) 
14'h2b69 : LOC =         127'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000010000000000000000000000; // D (0x00000000000000200000000000400000) 
14'h11c4 : LOC =         127'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000010000000000000000000000; // D (0x00000000000000400000000000400000) 
14'h27e9 : LOC =         127'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000010000000000000000000000; // D (0x00000000000000800000000000400000) 
14'h08c4 : LOC =         127'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000010000000000000000000000; // D (0x00000000000001000000000000400000) 
14'h15e9 : LOC =         127'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000010000000000000000000000; // D (0x00000000000002000000000000400000) 
14'h2fb3 : LOC =         127'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000010000000000000000000000; // D (0x00000000000004000000000000400000) 
14'h1870 : LOC =         127'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000010000000000000000000000; // D (0x00000000000008000000000000400000) 
14'h3481 : LOC =         127'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000010000000000000000000000; // D (0x00000000000010000000000000400000) 
14'h2e14 : LOC =         127'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000010000000000000000000000; // D (0x00000000000020000000000000400000) 
14'h1b3e : LOC =         127'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000010000000000000000000000; // D (0x00000000000040000000000000400000) 
14'h321d : LOC =         127'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000010000000000000000000000; // D (0x00000000000080000000000000400000) 
14'h232c : LOC =         127'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000010000000000000000000000; // D (0x00000000000100000000000000400000) 
14'h014e : LOC =         127'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000010000000000000000000000; // D (0x00000000000200000000000000400000) 
14'h06fd : LOC =         127'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000010000000000000000000000; // D (0x00000000000400000000000000400000) 
14'h099b : LOC =         127'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000010000000000000000000000; // D (0x00000000000800000000000000400000) 
14'h1757 : LOC =         127'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000010000000000000000000000; // D (0x00000000001000000000000000400000) 
14'h2acf : LOC =         127'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000010000000000000000000000; // D (0x00000000002000000000000000400000) 
14'h1288 : LOC =         127'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000010000000000000000000000; // D (0x00000000004000000000000000400000) 
14'h2171 : LOC =         127'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000010000000000000000000000; // D (0x00000000008000000000000000400000) 
14'h05f4 : LOC =         127'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000010000000000000000000000; // D (0x00000000010000000000000000400000) 
14'h0f89 : LOC =         127'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000010000000000000000000000; // D (0x00000000020000000000000000400000) 
14'h1b73 : LOC =         127'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000; // D (0x00000000040000000000000000400000) 
14'h3287 : LOC =         127'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000; // D (0x00000000080000000000000000400000) 
14'h2218 : LOC =         127'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000; // D (0x00000000100000000000000000400000) 
14'h0326 : LOC =         127'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000; // D (0x00000000200000000000000000400000) 
14'h022d : LOC =         127'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000; // D (0x00000000400000000000000000400000) 
14'h003b : LOC =         127'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000; // D (0x00000000800000000000000000400000) 
14'h0417 : LOC =         127'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000; // D (0x00000001000000000000000000400000) 
14'h0c4f : LOC =         127'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000; // D (0x00000002000000000000000000400000) 
14'h1cff : LOC =         127'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000; // D (0x00000004000000000000000000400000) 
14'h3d9f : LOC =         127'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000; // D (0x00000008000000000000000000400000) 
14'h3c28 : LOC =         127'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000; // D (0x00000010000000000000000000400000) 
14'h3f46 : LOC =         127'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000; // D (0x00000020000000000000000000400000) 
14'h399a : LOC =         127'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000; // D (0x00000040000000000000000000400000) 
14'h3422 : LOC =         127'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000; // D (0x00000080000000000000000000400000) 
14'h2f52 : LOC =         127'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000; // D (0x00000100000000000000000000400000) 
14'h19b2 : LOC =         127'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000; // D (0x00000200000000000000000000400000) 
14'h3705 : LOC =         127'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000; // D (0x00000400000000000000000000400000) 
14'h291c : LOC =         127'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000; // D (0x00000800000000000000000000400000) 
14'h152e : LOC =         127'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000; // D (0x00001000000000000000000000400000) 
14'h2e3d : LOC =         127'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000; // D (0x00002000000000000000000000400000) 
14'h1b6c : LOC =         127'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000; // D (0x00004000000000000000000000400000) 
14'h32b9 : LOC =         127'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000; // D (0x00008000000000000000000000400000) 
14'h2264 : LOC =         127'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000; // D (0x00010000000000000000000000400000) 
14'h03de : LOC =         127'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000; // D (0x00020000000000000000000000400000) 
14'h03dd : LOC =         127'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000; // D (0x00040000000000000000000000400000) 
14'h03db : LOC =         127'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000; // D (0x00080000000000000000000000400000) 
14'h03d7 : LOC =         127'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000; // D (0x00100000000000000000000000400000) 
14'h03cf : LOC =         127'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000; // D (0x00200000000000000000000000400000) 
14'h03ff : LOC =         127'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000; // D (0x00400000000000000000000000400000) 
14'h039f : LOC =         127'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000; // D (0x00800000000000000000000000400000) 
14'h035f : LOC =         127'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000; // D (0x01000000000000000000000000400000) 
14'h02df : LOC =         127'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000; // D (0x02000000000000000000000000400000) 
14'h01df : LOC =         127'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000; // D (0x04000000000000000000000000400000) 
14'h07df : LOC =         127'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000; // D (0x08000000000000000000000000400000) 
14'h0bdf : LOC =         127'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000; // D (0x10000000000000000000000000400000) 
14'h13df : LOC =         127'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000; // D (0x20000000000000000000000000400000) 
14'h23df : LOC =         127'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000; // D (0x40000000000000000000000000400000) 
14'h07be : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000; // S (0x00000000000000000000000000800000) 
14'h08c2 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000; // D (0x00000000000000000000000001800000) 
14'h1946 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000; // D (0x00000000000000000000000002800000) 
14'h3a4e : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000; // D (0x00000000000000000000000004800000) 
14'h3f29 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000100000000000000000000000; // D (0x00000000000000000000000008800000) 
14'h35e7 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000100000000000000000000000; // D (0x00000000000000000000000010800000) 
14'h207b : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000100000000000000000000000; // D (0x00000000000000000000000020800000) 
14'h0b43 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000100000000000000000000000; // D (0x00000000000000000000000040800000) 
14'h1e44 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000100000000000000000000000; // D (0x00000000000000000000000080800000) 
14'h344a : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000100000000000000000000000; // D (0x00000000000000000000000100800000) 
14'h2321 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000100000000000000000000000; // D (0x00000000000000000000000200800000) 
14'h0df7 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000100000000000000000000000; // D (0x00000000000000000000000400800000) 
14'h132c : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000100000000000000000000000; // D (0x00000000000000000000000800800000) 
14'h2e9a : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000100000000000000000000000; // D (0x00000000000000000000001000800000) 
14'h1681 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000100000000000000000000000; // D (0x00000000000000000000002000800000) 
14'h25c0 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000100000000000000000000000; // D (0x00000000000000000000004000800000) 
14'h0035 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000100000000000000000000000; // D (0x00000000000000000000008000800000) 
14'h08a8 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000100000000000000000000000; // D (0x00000000000000000000010000800000) 
14'h1992 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000100000000000000000000000; // D (0x00000000000000000000020000800000) 
14'h3be6 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000100000000000000000000000; // D (0x00000000000000000000040000800000) 
14'h3c79 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000100000000000000000000000; // D (0x00000000000000000000080000800000) 
14'h3347 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000100000000000000000000000; // D (0x00000000000000000000100000800000) 
14'h2d3b : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000100000000000000000000000; // D (0x00000000000000000000200000800000) 
14'h11c3 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000100000000000000000000000; // D (0x00000000000000000000400000800000) 
14'h2b44 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000100000000000000000000000; // D (0x00000000000000000000800000800000) 
14'h1d3d : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000100000000000000000000000; // D (0x00000000000000000001000000800000) 
14'h32b8 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000100000000000000000000000; // D (0x00000000000000000002000000800000) 
14'h2ec5 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000100000000000000000000000; // D (0x00000000000000000004000000800000) 
14'h163f : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000100000000000000000000000; // D (0x00000000000000000008000000800000) 
14'h24bc : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000100000000000000000000000; // D (0x00000000000000000010000000800000) 
14'h02cd : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000100000000000000000000000; // D (0x00000000000000000020000000800000) 
14'h0d58 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000100000000000000000000000; // D (0x00000000000000000040000000800000) 
14'h1272 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000100000000000000000000000; // D (0x00000000000000000080000000800000) 
14'h2c26 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000100000000000000000000000; // D (0x00000000000000000100000000800000) 
14'h13f9 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000100000000000000000000000; // D (0x00000000000000000200000000800000) 
14'h2f30 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000100000000000000000000000; // D (0x00000000000000000400000000800000) 
14'h15d5 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000100000000000000000000000; // D (0x00000000000000000800000000800000) 
14'h2368 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000100000000000000000000000; // D (0x00000000000000001000000000800000) 
14'h0d65 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000100000000000000000000000; // D (0x00000000000000002000000000800000) 
14'h1208 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000100000000000000000000000; // D (0x00000000000000004000000000800000) 
14'h2cd2 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000100000000000000000000000; // D (0x00000000000000008000000000800000) 
14'h1211 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000100000000000000000000000; // D (0x00000000000000010000000000800000) 
14'h2ce0 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000100000000000000000000000; // D (0x00000000000000020000000000800000) 
14'h1275 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000100000000000000000000000; // D (0x00000000000000040000000000800000) 
14'h2c28 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000100000000000000000000000; // D (0x00000000000000080000000000800000) 
14'h13e5 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000100000000000000000000000; // D (0x00000000000000100000000000800000) 
14'h2f08 : LOC =         127'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000100000000000000000000000; // D (0x00000000000000200000000000800000) 
14'h15a5 : LOC =         127'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000100000000000000000000000; // D (0x00000000000000400000000000800000) 
14'h2388 : LOC =         127'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000100000000000000000000000; // D (0x00000000000000800000000000800000) 
14'h0ca5 : LOC =         127'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000100000000000000000000000; // D (0x00000000000001000000000000800000) 
14'h1188 : LOC =         127'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000100000000000000000000000; // D (0x00000000000002000000000000800000) 
14'h2bd2 : LOC =         127'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000100000000000000000000000; // D (0x00000000000004000000000000800000) 
14'h1c11 : LOC =         127'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000100000000000000000000000; // D (0x00000000000008000000000000800000) 
14'h30e0 : LOC =         127'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000100000000000000000000000; // D (0x00000000000010000000000000800000) 
14'h2a75 : LOC =         127'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000100000000000000000000000; // D (0x00000000000020000000000000800000) 
14'h1f5f : LOC =         127'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000100000000000000000000000; // D (0x00000000000040000000000000800000) 
14'h367c : LOC =         127'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000100000000000000000000000; // D (0x00000000000080000000000000800000) 
14'h274d : LOC =         127'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000100000000000000000000000; // D (0x00000000000100000000000000800000) 
14'h052f : LOC =         127'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000100000000000000000000000; // D (0x00000000000200000000000000800000) 
14'h029c : LOC =         127'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000100000000000000000000000; // D (0x00000000000400000000000000800000) 
14'h0dfa : LOC =         127'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000100000000000000000000000; // D (0x00000000000800000000000000800000) 
14'h1336 : LOC =         127'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000100000000000000000000000; // D (0x00000000001000000000000000800000) 
14'h2eae : LOC =         127'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000100000000000000000000000; // D (0x00000000002000000000000000800000) 
14'h16e9 : LOC =         127'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000100000000000000000000000; // D (0x00000000004000000000000000800000) 
14'h2510 : LOC =         127'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000100000000000000000000000; // D (0x00000000008000000000000000800000) 
14'h0195 : LOC =         127'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000100000000000000000000000; // D (0x00000000010000000000000000800000) 
14'h0be8 : LOC =         127'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000100000000000000000000000; // D (0x00000000020000000000000000800000) 
14'h1f12 : LOC =         127'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000; // D (0x00000000040000000000000000800000) 
14'h36e6 : LOC =         127'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000; // D (0x00000000080000000000000000800000) 
14'h2679 : LOC =         127'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000; // D (0x00000000100000000000000000800000) 
14'h0747 : LOC =         127'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000; // D (0x00000000200000000000000000800000) 
14'h064c : LOC =         127'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000; // D (0x00000000400000000000000000800000) 
14'h045a : LOC =         127'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000; // D (0x00000000800000000000000000800000) 
14'h0076 : LOC =         127'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000; // D (0x00000001000000000000000000800000) 
14'h082e : LOC =         127'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000; // D (0x00000002000000000000000000800000) 
14'h189e : LOC =         127'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000; // D (0x00000004000000000000000000800000) 
14'h39fe : LOC =         127'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000; // D (0x00000008000000000000000000800000) 
14'h3849 : LOC =         127'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000; // D (0x00000010000000000000000000800000) 
14'h3b27 : LOC =         127'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000; // D (0x00000020000000000000000000800000) 
14'h3dfb : LOC =         127'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000; // D (0x00000040000000000000000000800000) 
14'h3043 : LOC =         127'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000; // D (0x00000080000000000000000000800000) 
14'h2b33 : LOC =         127'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000; // D (0x00000100000000000000000000800000) 
14'h1dd3 : LOC =         127'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000; // D (0x00000200000000000000000000800000) 
14'h3364 : LOC =         127'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000; // D (0x00000400000000000000000000800000) 
14'h2d7d : LOC =         127'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000; // D (0x00000800000000000000000000800000) 
14'h114f : LOC =         127'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000; // D (0x00001000000000000000000000800000) 
14'h2a5c : LOC =         127'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000; // D (0x00002000000000000000000000800000) 
14'h1f0d : LOC =         127'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000; // D (0x00004000000000000000000000800000) 
14'h36d8 : LOC =         127'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000; // D (0x00008000000000000000000000800000) 
14'h2605 : LOC =         127'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000; // D (0x00010000000000000000000000800000) 
14'h07bf : LOC =         127'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000; // D (0x00020000000000000000000000800000) 
14'h07bc : LOC =         127'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000; // D (0x00040000000000000000000000800000) 
14'h07ba : LOC =         127'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000; // D (0x00080000000000000000000000800000) 
14'h07b6 : LOC =         127'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000; // D (0x00100000000000000000000000800000) 
14'h07ae : LOC =         127'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000; // D (0x00200000000000000000000000800000) 
14'h079e : LOC =         127'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000; // D (0x00400000000000000000000000800000) 
14'h07fe : LOC =         127'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000; // D (0x00800000000000000000000000800000) 
14'h073e : LOC =         127'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000; // D (0x01000000000000000000000000800000) 
14'h06be : LOC =         127'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000; // D (0x02000000000000000000000000800000) 
14'h05be : LOC =         127'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000; // D (0x04000000000000000000000000800000) 
14'h03be : LOC =         127'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000; // D (0x08000000000000000000000000800000) 
14'h0fbe : LOC =         127'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000; // D (0x10000000000000000000000000800000) 
14'h17be : LOC =         127'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000; // D (0x20000000000000000000000000800000) 
14'h27be : LOC =         127'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000; // D (0x40000000000000000000000000800000) 
14'h0f7c : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000; // S (0x00000000000000000000000001000000) 
14'h1184 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000; // D (0x00000000000000000000000003000000) 
14'h328c : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000000000000000000000000; // D (0x00000000000000000000000005000000) 
14'h37eb : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000000000; // D (0x00000000000000000000000009000000) 
14'h3d25 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000000000000000000000000; // D (0x00000000000000000000000011000000) 
14'h28b9 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100001000000000000000000000000; // D (0x00000000000000000000000021000000) 
14'h0381 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000001000000000000000000000000; // D (0x00000000000000000000000041000000) 
14'h1686 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000001000000000000000000000000; // D (0x00000000000000000000000081000000) 
14'h3c88 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000001000000000000000000000000; // D (0x00000000000000000000000101000000) 
14'h2be3 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000001000000000000000000000000; // D (0x00000000000000000000000201000000) 
14'h0535 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000001000000000000000000000000; // D (0x00000000000000000000000401000000) 
14'h1bee : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000001000000000000000000000000; // D (0x00000000000000000000000801000000) 
14'h2658 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000001000000000000000000000000; // D (0x00000000000000000000001001000000) 
14'h1e43 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000001000000000000000000000000; // D (0x00000000000000000000002001000000) 
14'h2d02 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000001000000000000000000000000; // D (0x00000000000000000000004001000000) 
14'h08f7 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000001000000000000000000000000; // D (0x00000000000000000000008001000000) 
14'h006a : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001000000000000000000000000; // D (0x00000000000000000000010001000000) 
14'h1150 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000001000000000000000000000000; // D (0x00000000000000000000020001000000) 
14'h3324 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000001000000000000000000000000; // D (0x00000000000000000000040001000000) 
14'h34bb : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000001000000000000000000000000; // D (0x00000000000000000000080001000000) 
14'h3b85 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000001000000000000000000000000; // D (0x00000000000000000000100001000000) 
14'h25f9 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000001000000000000000000000000; // D (0x00000000000000000000200001000000) 
14'h1901 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000001000000000000000000000000; // D (0x00000000000000000000400001000000) 
14'h2386 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000001000000000000000000000000; // D (0x00000000000000000000800001000000) 
14'h15ff : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000001000000000000000000000000; // D (0x00000000000000000001000001000000) 
14'h3a7a : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000001000000000000000000000000; // D (0x00000000000000000002000001000000) 
14'h2607 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000001000000000000000000000000; // D (0x00000000000000000004000001000000) 
14'h1efd : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000001000000000000000000000000; // D (0x00000000000000000008000001000000) 
14'h2c7e : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000001000000000000000000000000; // D (0x00000000000000000010000001000000) 
14'h0a0f : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000001000000000000000000000000; // D (0x00000000000000000020000001000000) 
14'h059a : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000001000000000000000000000000; // D (0x00000000000000000040000001000000) 
14'h1ab0 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000001000000000000000000000000; // D (0x00000000000000000080000001000000) 
14'h24e4 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000001000000000000000000000000; // D (0x00000000000000000100000001000000) 
14'h1b3b : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000001000000000000000000000000; // D (0x00000000000000000200000001000000) 
14'h27f2 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000001000000000000000000000000; // D (0x00000000000000000400000001000000) 
14'h1d17 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000001000000000000000000000000; // D (0x00000000000000000800000001000000) 
14'h2baa : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000001000000000000000000000000; // D (0x00000000000000001000000001000000) 
14'h05a7 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000001000000000000000000000000; // D (0x00000000000000002000000001000000) 
14'h1aca : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000000000000000000; // D (0x00000000000000004000000001000000) 
14'h2410 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000001000000000000000000000000; // D (0x00000000000000008000000001000000) 
14'h1ad3 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000001000000000000000000000000; // D (0x00000000000000010000000001000000) 
14'h2422 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000001000000000000000000000000; // D (0x00000000000000020000000001000000) 
14'h1ab7 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000001000000000000000000000000; // D (0x00000000000000040000000001000000) 
14'h24ea : LOC =         127'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000001000000000000000000000000; // D (0x00000000000000080000000001000000) 
14'h1b27 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000001000000000000000000000000; // D (0x00000000000000100000000001000000) 
14'h27ca : LOC =         127'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000001000000000000000000000000; // D (0x00000000000000200000000001000000) 
14'h1d67 : LOC =         127'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000001000000000000000000000000; // D (0x00000000000000400000000001000000) 
14'h2b4a : LOC =         127'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000001000000000000000000000000; // D (0x00000000000000800000000001000000) 
14'h0467 : LOC =         127'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000001000000000000000000000000; // D (0x00000000000001000000000001000000) 
14'h194a : LOC =         127'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000001000000000000000000000000; // D (0x00000000000002000000000001000000) 
14'h2310 : LOC =         127'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000001000000000000000000000000; // D (0x00000000000004000000000001000000) 
14'h14d3 : LOC =         127'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000001000000000000000000000000; // D (0x00000000000008000000000001000000) 
14'h3822 : LOC =         127'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000001000000000000000000000000; // D (0x00000000000010000000000001000000) 
14'h22b7 : LOC =         127'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000001000000000000000000000000; // D (0x00000000000020000000000001000000) 
14'h179d : LOC =         127'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000001000000000000000000000000; // D (0x00000000000040000000000001000000) 
14'h3ebe : LOC =         127'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000001000000000000000000000000; // D (0x00000000000080000000000001000000) 
14'h2f8f : LOC =         127'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000001000000000000000000000000; // D (0x00000000000100000000000001000000) 
14'h0ded : LOC =         127'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000001000000000000000000000000; // D (0x00000000000200000000000001000000) 
14'h0a5e : LOC =         127'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000001000000000000000000000000; // D (0x00000000000400000000000001000000) 
14'h0538 : LOC =         127'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000001000000000000000000000000; // D (0x00000000000800000000000001000000) 
14'h1bf4 : LOC =         127'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000001000000000000000000000000; // D (0x00000000001000000000000001000000) 
14'h266c : LOC =         127'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000001000000000000000000000000; // D (0x00000000002000000000000001000000) 
14'h1e2b : LOC =         127'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000001000000000000000000000000; // D (0x00000000004000000000000001000000) 
14'h2dd2 : LOC =         127'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000001000000000000000000000000; // D (0x00000000008000000000000001000000) 
14'h0957 : LOC =         127'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000001000000000000000000000000; // D (0x00000000010000000000000001000000) 
14'h032a : LOC =         127'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000001000000000000000000000000; // D (0x00000000020000000000000001000000) 
14'h17d0 : LOC =         127'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000; // D (0x00000000040000000000000001000000) 
14'h3e24 : LOC =         127'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000; // D (0x00000000080000000000000001000000) 
14'h2ebb : LOC =         127'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000; // D (0x00000000100000000000000001000000) 
14'h0f85 : LOC =         127'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000; // D (0x00000000200000000000000001000000) 
14'h0e8e : LOC =         127'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000; // D (0x00000000400000000000000001000000) 
14'h0c98 : LOC =         127'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000; // D (0x00000000800000000000000001000000) 
14'h08b4 : LOC =         127'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000; // D (0x00000001000000000000000001000000) 
14'h00ec : LOC =         127'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000; // D (0x00000002000000000000000001000000) 
14'h105c : LOC =         127'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000; // D (0x00000004000000000000000001000000) 
14'h313c : LOC =         127'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000; // D (0x00000008000000000000000001000000) 
14'h308b : LOC =         127'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000; // D (0x00000010000000000000000001000000) 
14'h33e5 : LOC =         127'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000; // D (0x00000020000000000000000001000000) 
14'h3539 : LOC =         127'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000; // D (0x00000040000000000000000001000000) 
14'h3881 : LOC =         127'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000; // D (0x00000080000000000000000001000000) 
14'h23f1 : LOC =         127'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000; // D (0x00000100000000000000000001000000) 
14'h1511 : LOC =         127'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000; // D (0x00000200000000000000000001000000) 
14'h3ba6 : LOC =         127'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000; // D (0x00000400000000000000000001000000) 
14'h25bf : LOC =         127'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000; // D (0x00000800000000000000000001000000) 
14'h198d : LOC =         127'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000; // D (0x00001000000000000000000001000000) 
14'h229e : LOC =         127'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000; // D (0x00002000000000000000000001000000) 
14'h17cf : LOC =         127'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000; // D (0x00004000000000000000000001000000) 
14'h3e1a : LOC =         127'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000; // D (0x00008000000000000000000001000000) 
14'h2ec7 : LOC =         127'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000; // D (0x00010000000000000000000001000000) 
14'h0f7d : LOC =         127'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000; // D (0x00020000000000000000000001000000) 
14'h0f7e : LOC =         127'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000; // D (0x00040000000000000000000001000000) 
14'h0f78 : LOC =         127'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000; // D (0x00080000000000000000000001000000) 
14'h0f74 : LOC =         127'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000; // D (0x00100000000000000000000001000000) 
14'h0f6c : LOC =         127'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000; // D (0x00200000000000000000000001000000) 
14'h0f5c : LOC =         127'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000; // D (0x00400000000000000000000001000000) 
14'h0f3c : LOC =         127'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000; // D (0x00800000000000000000000001000000) 
14'h0ffc : LOC =         127'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000; // D (0x01000000000000000000000001000000) 
14'h0e7c : LOC =         127'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000; // D (0x02000000000000000000000001000000) 
14'h0d7c : LOC =         127'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000; // D (0x04000000000000000000000001000000) 
14'h0b7c : LOC =         127'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000; // D (0x08000000000000000000000001000000) 
14'h077c : LOC =         127'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000; // D (0x10000000000000000000000001000000) 
14'h1f7c : LOC =         127'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000; // D (0x20000000000000000000000001000000) 
14'h2f7c : LOC =         127'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000; // D (0x40000000000000000000000001000000) 
14'h1ef8 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000; // S (0x00000000000000000000000002000000) 
14'h2308 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000000; // D (0x00000000000000000000000006000000) 
14'h266f : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000000000000000000000000; // D (0x0000000000000000000000000a000000) 
14'h2ca1 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000; // D (0x00000000000000000000000012000000) 
14'h393d : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010000000000000000000000000; // D (0x00000000000000000000000022000000) 
14'h1205 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000010000000000000000000000000; // D (0x00000000000000000000000042000000) 
14'h0702 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000010000000000000000000000000; // D (0x00000000000000000000000082000000) 
14'h2d0c : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000010000000000000000000000000; // D (0x00000000000000000000000102000000) 
14'h3a67 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000010000000000000000000000000; // D (0x00000000000000000000000202000000) 
14'h14b1 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000010000000000000000000000000; // D (0x00000000000000000000000402000000) 
14'h0a6a : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000010000000000000000000000000; // D (0x00000000000000000000000802000000) 
14'h37dc : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000010000000000000000000000000; // D (0x00000000000000000000001002000000) 
14'h0fc7 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000010000000000000000000000000; // D (0x00000000000000000000002002000000) 
14'h3c86 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000010000000000000000000000000; // D (0x00000000000000000000004002000000) 
14'h1973 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000010000000000000000000000000; // D (0x00000000000000000000008002000000) 
14'h11ee : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000010000000000000000000000000; // D (0x00000000000000000000010002000000) 
14'h00d4 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000010000000000000000000000000; // D (0x00000000000000000000020002000000) 
14'h22a0 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000010000000000000000000000000; // D (0x00000000000000000000040002000000) 
14'h253f : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000010000000000000000000000000; // D (0x00000000000000000000080002000000) 
14'h2a01 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000010000000000000000000000000; // D (0x00000000000000000000100002000000) 
14'h347d : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000010000000000000000000000000; // D (0x00000000000000000000200002000000) 
14'h0885 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000010000000000000000000000000; // D (0x00000000000000000000400002000000) 
14'h3202 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000010000000000000000000000000; // D (0x00000000000000000000800002000000) 
14'h047b : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000010000000000000000000000000; // D (0x00000000000000000001000002000000) 
14'h2bfe : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000010000000000000000000000000; // D (0x00000000000000000002000002000000) 
14'h3783 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000010000000000000000000000000; // D (0x00000000000000000004000002000000) 
14'h0f79 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000010000000000000000000000000; // D (0x00000000000000000008000002000000) 
14'h3dfa : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000010000000000000000000000000; // D (0x00000000000000000010000002000000) 
14'h1b8b : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000010000000000000000000000000; // D (0x00000000000000000020000002000000) 
14'h141e : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000010000000000000000000000000; // D (0x00000000000000000040000002000000) 
14'h0b34 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000010000000000000000000000000; // D (0x00000000000000000080000002000000) 
14'h3560 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000010000000000000000000000000; // D (0x00000000000000000100000002000000) 
14'h0abf : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000010000000000000000000000000; // D (0x00000000000000000200000002000000) 
14'h3676 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000010000000000000000000000000; // D (0x00000000000000000400000002000000) 
14'h0c93 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000; // D (0x00000000000000000800000002000000) 
14'h3a2e : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000010000000000000000000000000; // D (0x00000000000000001000000002000000) 
14'h1423 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000010000000000000000000000000; // D (0x00000000000000002000000002000000) 
14'h0b4e : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000; // D (0x00000000000000004000000002000000) 
14'h3594 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000010000000000000000000000000; // D (0x00000000000000008000000002000000) 
14'h0b57 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000010000000000000000000000000; // D (0x00000000000000010000000002000000) 
14'h35a6 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000010000000000000000000000000; // D (0x00000000000000020000000002000000) 
14'h0b33 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000010000000000000000000000000; // D (0x00000000000000040000000002000000) 
14'h356e : LOC =         127'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000010000000000000000000000000; // D (0x00000000000000080000000002000000) 
14'h0aa3 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000010000000000000000000000000; // D (0x00000000000000100000000002000000) 
14'h364e : LOC =         127'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000010000000000000000000000000; // D (0x00000000000000200000000002000000) 
14'h0ce3 : LOC =         127'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000010000000000000000000000000; // D (0x00000000000000400000000002000000) 
14'h3ace : LOC =         127'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000010000000000000000000000000; // D (0x00000000000000800000000002000000) 
14'h15e3 : LOC =         127'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000010000000000000000000000000; // D (0x00000000000001000000000002000000) 
14'h08ce : LOC =         127'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000010000000000000000000000000; // D (0x00000000000002000000000002000000) 
14'h3294 : LOC =         127'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000010000000000000000000000000; // D (0x00000000000004000000000002000000) 
14'h0557 : LOC =         127'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000010000000000000000000000000; // D (0x00000000000008000000000002000000) 
14'h29a6 : LOC =         127'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000010000000000000000000000000; // D (0x00000000000010000000000002000000) 
14'h3333 : LOC =         127'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000010000000000000000000000000; // D (0x00000000000020000000000002000000) 
14'h0619 : LOC =         127'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000010000000000000000000000000; // D (0x00000000000040000000000002000000) 
14'h2f3a : LOC =         127'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000010000000000000000000000000; // D (0x00000000000080000000000002000000) 
14'h3e0b : LOC =         127'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000010000000000000000000000000; // D (0x00000000000100000000000002000000) 
14'h1c69 : LOC =         127'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000010000000000000000000000000; // D (0x00000000000200000000000002000000) 
14'h1bda : LOC =         127'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000010000000000000000000000000; // D (0x00000000000400000000000002000000) 
14'h14bc : LOC =         127'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000010000000000000000000000000; // D (0x00000000000800000000000002000000) 
14'h0a70 : LOC =         127'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000010000000000000000000000000; // D (0x00000000001000000000000002000000) 
14'h37e8 : LOC =         127'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000010000000000000000000000000; // D (0x00000000002000000000000002000000) 
14'h0faf : LOC =         127'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000010000000000000000000000000; // D (0x00000000004000000000000002000000) 
14'h3c56 : LOC =         127'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000010000000000000000000000000; // D (0x00000000008000000000000002000000) 
14'h18d3 : LOC =         127'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000010000000000000000000000000; // D (0x00000000010000000000000002000000) 
14'h12ae : LOC =         127'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000010000000000000000000000000; // D (0x00000000020000000000000002000000) 
14'h0654 : LOC =         127'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000; // D (0x00000000040000000000000002000000) 
14'h2fa0 : LOC =         127'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000; // D (0x00000000080000000000000002000000) 
14'h3f3f : LOC =         127'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000; // D (0x00000000100000000000000002000000) 
14'h1e01 : LOC =         127'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000; // D (0x00000000200000000000000002000000) 
14'h1f0a : LOC =         127'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000; // D (0x00000000400000000000000002000000) 
14'h1d1c : LOC =         127'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000; // D (0x00000000800000000000000002000000) 
14'h1930 : LOC =         127'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000; // D (0x00000001000000000000000002000000) 
14'h1168 : LOC =         127'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000; // D (0x00000002000000000000000002000000) 
14'h01d8 : LOC =         127'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000; // D (0x00000004000000000000000002000000) 
14'h20b8 : LOC =         127'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000; // D (0x00000008000000000000000002000000) 
14'h210f : LOC =         127'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000; // D (0x00000010000000000000000002000000) 
14'h2261 : LOC =         127'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000; // D (0x00000020000000000000000002000000) 
14'h24bd : LOC =         127'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000; // D (0x00000040000000000000000002000000) 
14'h2905 : LOC =         127'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000; // D (0x00000080000000000000000002000000) 
14'h3275 : LOC =         127'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000; // D (0x00000100000000000000000002000000) 
14'h0495 : LOC =         127'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000; // D (0x00000200000000000000000002000000) 
14'h2a22 : LOC =         127'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000; // D (0x00000400000000000000000002000000) 
14'h343b : LOC =         127'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000; // D (0x00000800000000000000000002000000) 
14'h0809 : LOC =         127'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000; // D (0x00001000000000000000000002000000) 
14'h331a : LOC =         127'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000; // D (0x00002000000000000000000002000000) 
14'h064b : LOC =         127'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000; // D (0x00004000000000000000000002000000) 
14'h2f9e : LOC =         127'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000; // D (0x00008000000000000000000002000000) 
14'h3f43 : LOC =         127'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000; // D (0x00010000000000000000000002000000) 
14'h1ef9 : LOC =         127'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000; // D (0x00020000000000000000000002000000) 
14'h1efa : LOC =         127'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000; // D (0x00040000000000000000000002000000) 
14'h1efc : LOC =         127'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000; // D (0x00080000000000000000000002000000) 
14'h1ef0 : LOC =         127'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000; // D (0x00100000000000000000000002000000) 
14'h1ee8 : LOC =         127'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000; // D (0x00200000000000000000000002000000) 
14'h1ed8 : LOC =         127'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000; // D (0x00400000000000000000000002000000) 
14'h1eb8 : LOC =         127'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000; // D (0x00800000000000000000000002000000) 
14'h1e78 : LOC =         127'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000; // D (0x01000000000000000000000002000000) 
14'h1ff8 : LOC =         127'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000; // D (0x02000000000000000000000002000000) 
14'h1cf8 : LOC =         127'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000; // D (0x04000000000000000000000002000000) 
14'h1af8 : LOC =         127'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000; // D (0x08000000000000000000000002000000) 
14'h16f8 : LOC =         127'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000; // D (0x10000000000000000000000002000000) 
14'h0ef8 : LOC =         127'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000; // D (0x20000000000000000000000002000000) 
14'h3ef8 : LOC =         127'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000; // D (0x40000000000000000000000002000000) 
14'h3df0 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000; // S (0x00000000000000000000000004000000) 
14'h0567 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000; // D (0x0000000000000000000000000c000000) 
14'h0fa9 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000; // D (0x00000000000000000000000014000000) 
14'h1a35 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000; // D (0x00000000000000000000000024000000) 
14'h310d : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000100000000000000000000000000; // D (0x00000000000000000000000044000000) 
14'h240a : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000100000000000000000000000000; // D (0x00000000000000000000000084000000) 
14'h0e04 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000100000000000000000000000000; // D (0x00000000000000000000000104000000) 
14'h196f : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000100000000000000000000000000; // D (0x00000000000000000000000204000000) 
14'h37b9 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000100000000000000000000000000; // D (0x00000000000000000000000404000000) 
14'h2962 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000100000000000000000000000000; // D (0x00000000000000000000000804000000) 
14'h14d4 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000100000000000000000000000000; // D (0x00000000000000000000001004000000) 
14'h2ccf : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000100000000000000000000000000; // D (0x00000000000000000000002004000000) 
14'h1f8e : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000100000000000000000000000000; // D (0x00000000000000000000004004000000) 
14'h3a7b : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000100000000000000000000000000; // D (0x00000000000000000000008004000000) 
14'h32e6 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000100000000000000000000000000; // D (0x00000000000000000000010004000000) 
14'h23dc : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000100000000000000000000000000; // D (0x00000000000000000000020004000000) 
14'h01a8 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000100000000000000000000000000; // D (0x00000000000000000000040004000000) 
14'h0637 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000100000000000000000000000000; // D (0x00000000000000000000080004000000) 
14'h0909 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000100000000000000000000000000; // D (0x00000000000000000000100004000000) 
14'h1775 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000100000000000000000000000000; // D (0x00000000000000000000200004000000) 
14'h2b8d : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000100000000000000000000000000; // D (0x00000000000000000000400004000000) 
14'h110a : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000100000000000000000000000000; // D (0x00000000000000000000800004000000) 
14'h2773 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000100000000000000000000000000; // D (0x00000000000000000001000004000000) 
14'h08f6 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000100000000000000000000000000; // D (0x00000000000000000002000004000000) 
14'h148b : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000100000000000000000000000000; // D (0x00000000000000000004000004000000) 
14'h2c71 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000100000000000000000000000000; // D (0x00000000000000000008000004000000) 
14'h1ef2 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000100000000000000000000000000; // D (0x00000000000000000010000004000000) 
14'h3883 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000100000000000000000000000000; // D (0x00000000000000000020000004000000) 
14'h3716 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000100000000000000000000000000; // D (0x00000000000000000040000004000000) 
14'h283c : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000100000000000000000000000000; // D (0x00000000000000000080000004000000) 
14'h1668 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000100000000000000000000000000; // D (0x00000000000000000100000004000000) 
14'h29b7 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000100000000000000000000000000; // D (0x00000000000000000200000004000000) 
14'h157e : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000100000000000000000000000000; // D (0x00000000000000000400000004000000) 
14'h2f9b : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000100000000000000000000000000; // D (0x00000000000000000800000004000000) 
14'h1926 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000100000000000000000000000000; // D (0x00000000000000001000000004000000) 
14'h372b : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000100000000000000000000000000; // D (0x00000000000000002000000004000000) 
14'h2846 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000100000000000000000000000000; // D (0x00000000000000004000000004000000) 
14'h169c : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000100000000000000000000000000; // D (0x00000000000000008000000004000000) 
14'h285f : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000100000000000000000000000000; // D (0x00000000000000010000000004000000) 
14'h16ae : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000100000000000000000000000000; // D (0x00000000000000020000000004000000) 
14'h283b : LOC =         127'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000100000000000000000000000000; // D (0x00000000000000040000000004000000) 
14'h1666 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000100000000000000000000000000; // D (0x00000000000000080000000004000000) 
14'h29ab : LOC =         127'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000100000000000000000000000000; // D (0x00000000000000100000000004000000) 
14'h1546 : LOC =         127'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000100000000000000000000000000; // D (0x00000000000000200000000004000000) 
14'h2feb : LOC =         127'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000100000000000000000000000000; // D (0x00000000000000400000000004000000) 
14'h19c6 : LOC =         127'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000100000000000000000000000000; // D (0x00000000000000800000000004000000) 
14'h36eb : LOC =         127'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000100000000000000000000000000; // D (0x00000000000001000000000004000000) 
14'h2bc6 : LOC =         127'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000100000000000000000000000000; // D (0x00000000000002000000000004000000) 
14'h119c : LOC =         127'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000100000000000000000000000000; // D (0x00000000000004000000000004000000) 
14'h265f : LOC =         127'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000100000000000000000000000000; // D (0x00000000000008000000000004000000) 
14'h0aae : LOC =         127'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000100000000000000000000000000; // D (0x00000000000010000000000004000000) 
14'h103b : LOC =         127'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000100000000000000000000000000; // D (0x00000000000020000000000004000000) 
14'h2511 : LOC =         127'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000100000000000000000000000000; // D (0x00000000000040000000000004000000) 
14'h0c32 : LOC =         127'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000100000000000000000000000000; // D (0x00000000000080000000000004000000) 
14'h1d03 : LOC =         127'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000100000000000000000000000000; // D (0x00000000000100000000000004000000) 
14'h3f61 : LOC =         127'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000100000000000000000000000000; // D (0x00000000000200000000000004000000) 
14'h38d2 : LOC =         127'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000100000000000000000000000000; // D (0x00000000000400000000000004000000) 
14'h37b4 : LOC =         127'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000100000000000000000000000000; // D (0x00000000000800000000000004000000) 
14'h2978 : LOC =         127'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000100000000000000000000000000; // D (0x00000000001000000000000004000000) 
14'h14e0 : LOC =         127'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000100000000000000000000000000; // D (0x00000000002000000000000004000000) 
14'h2ca7 : LOC =         127'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000100000000000000000000000000; // D (0x00000000004000000000000004000000) 
14'h1f5e : LOC =         127'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000100000000000000000000000000; // D (0x00000000008000000000000004000000) 
14'h3bdb : LOC =         127'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000100000000000000000000000000; // D (0x00000000010000000000000004000000) 
14'h31a6 : LOC =         127'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000100000000000000000000000000; // D (0x00000000020000000000000004000000) 
14'h255c : LOC =         127'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000; // D (0x00000000040000000000000004000000) 
14'h0ca8 : LOC =         127'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000; // D (0x00000000080000000000000004000000) 
14'h1c37 : LOC =         127'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000; // D (0x00000000100000000000000004000000) 
14'h3d09 : LOC =         127'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000; // D (0x00000000200000000000000004000000) 
14'h3c02 : LOC =         127'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000; // D (0x00000000400000000000000004000000) 
14'h3e14 : LOC =         127'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000; // D (0x00000000800000000000000004000000) 
14'h3a38 : LOC =         127'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000; // D (0x00000001000000000000000004000000) 
14'h3260 : LOC =         127'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000; // D (0x00000002000000000000000004000000) 
14'h22d0 : LOC =         127'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000; // D (0x00000004000000000000000004000000) 
14'h03b0 : LOC =         127'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000; // D (0x00000008000000000000000004000000) 
14'h0207 : LOC =         127'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000; // D (0x00000010000000000000000004000000) 
14'h0169 : LOC =         127'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000; // D (0x00000020000000000000000004000000) 
14'h07b5 : LOC =         127'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000; // D (0x00000040000000000000000004000000) 
14'h0a0d : LOC =         127'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000; // D (0x00000080000000000000000004000000) 
14'h117d : LOC =         127'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000; // D (0x00000100000000000000000004000000) 
14'h279d : LOC =         127'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000; // D (0x00000200000000000000000004000000) 
14'h092a : LOC =         127'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000; // D (0x00000400000000000000000004000000) 
14'h1733 : LOC =         127'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000; // D (0x00000800000000000000000004000000) 
14'h2b01 : LOC =         127'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000; // D (0x00001000000000000000000004000000) 
14'h1012 : LOC =         127'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000; // D (0x00002000000000000000000004000000) 
14'h2543 : LOC =         127'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000; // D (0x00004000000000000000000004000000) 
14'h0c96 : LOC =         127'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000; // D (0x00008000000000000000000004000000) 
14'h1c4b : LOC =         127'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000; // D (0x00010000000000000000000004000000) 
14'h3df1 : LOC =         127'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000; // D (0x00020000000000000000000004000000) 
14'h3df2 : LOC =         127'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000; // D (0x00040000000000000000000004000000) 
14'h3df4 : LOC =         127'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000; // D (0x00080000000000000000000004000000) 
14'h3df8 : LOC =         127'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000; // D (0x00100000000000000000000004000000) 
14'h3de0 : LOC =         127'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000; // D (0x00200000000000000000000004000000) 
14'h3dd0 : LOC =         127'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000; // D (0x00400000000000000000000004000000) 
14'h3db0 : LOC =         127'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000; // D (0x00800000000000000000000004000000) 
14'h3d70 : LOC =         127'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000; // D (0x01000000000000000000000004000000) 
14'h3cf0 : LOC =         127'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000; // D (0x02000000000000000000000004000000) 
14'h3ff0 : LOC =         127'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000; // D (0x04000000000000000000000004000000) 
14'h39f0 : LOC =         127'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000; // D (0x08000000000000000000000004000000) 
14'h35f0 : LOC =         127'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000; // D (0x10000000000000000000000004000000) 
14'h2df0 : LOC =         127'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000; // D (0x20000000000000000000000004000000) 
14'h1df0 : LOC =         127'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000; // D (0x40000000000000000000000004000000) 
14'h3897 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000; // S (0x00000000000000000000000008000000) 
14'h0ace : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000000; // D (0x00000000000000000000000018000000) 
14'h1f52 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000000000000000000000000000; // D (0x00000000000000000000000028000000) 
14'h346a : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000; // D (0x00000000000000000000000048000000) 
14'h216d : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000000000000000000000000000; // D (0x00000000000000000000000088000000) 
14'h0b63 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100001000000000000000000000000000; // D (0x00000000000000000000000108000000) 
14'h1c08 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000001000000000000000000000000000; // D (0x00000000000000000000000208000000) 
14'h32de : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000001000000000000000000000000000; // D (0x00000000000000000000000408000000) 
14'h2c05 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000001000000000000000000000000000; // D (0x00000000000000000000000808000000) 
14'h11b3 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000001000000000000000000000000000; // D (0x00000000000000000000001008000000) 
14'h29a8 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000001000000000000000000000000000; // D (0x00000000000000000000002008000000) 
14'h1ae9 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000001000000000000000000000000000; // D (0x00000000000000000000004008000000) 
14'h3f1c : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000001000000000000000000000000000; // D (0x00000000000000000000008008000000) 
14'h3781 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000001000000000000000000000000000; // D (0x00000000000000000000010008000000) 
14'h26bb : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000001000000000000000000000000000; // D (0x00000000000000000000020008000000) 
14'h04cf : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000001000000000000000000000000000; // D (0x00000000000000000000040008000000) 
14'h0350 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001000000000000000000000000000; // D (0x00000000000000000000080008000000) 
14'h0c6e : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000001000000000000000000000000000; // D (0x00000000000000000000100008000000) 
14'h1212 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000001000000000000000000000000000; // D (0x00000000000000000000200008000000) 
14'h2eea : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000001000000000000000000000000000; // D (0x00000000000000000000400008000000) 
14'h146d : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000001000000000000000000000000000; // D (0x00000000000000000000800008000000) 
14'h2214 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000001000000000000000000000000000; // D (0x00000000000000000001000008000000) 
14'h0d91 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000001000000000000000000000000000; // D (0x00000000000000000002000008000000) 
14'h11ec : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000001000000000000000000000000000; // D (0x00000000000000000004000008000000) 
14'h2916 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000001000000000000000000000000000; // D (0x00000000000000000008000008000000) 
14'h1b95 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000001000000000000000000000000000; // D (0x00000000000000000010000008000000) 
14'h3de4 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000001000000000000000000000000000; // D (0x00000000000000000020000008000000) 
14'h3271 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000001000000000000000000000000000; // D (0x00000000000000000040000008000000) 
14'h2d5b : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000001000000000000000000000000000; // D (0x00000000000000000080000008000000) 
14'h130f : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000001000000000000000000000000000; // D (0x00000000000000000100000008000000) 
14'h2cd0 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000001000000000000000000000000000; // D (0x00000000000000000200000008000000) 
14'h1019 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000001000000000000000000000000000; // D (0x00000000000000000400000008000000) 
14'h2afc : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000001000000000000000000000000000; // D (0x00000000000000000800000008000000) 
14'h1c41 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000001000000000000000000000000000; // D (0x00000000000000001000000008000000) 
14'h324c : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000001000000000000000000000000000; // D (0x00000000000000002000000008000000) 
14'h2d21 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000001000000000000000000000000000; // D (0x00000000000000004000000008000000) 
14'h13fb : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000001000000000000000000000000000; // D (0x00000000000000008000000008000000) 
14'h2d38 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000001000000000000000000000000000; // D (0x00000000000000010000000008000000) 
14'h13c9 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000000000000000000000; // D (0x00000000000000020000000008000000) 
14'h2d5c : LOC =         127'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000001000000000000000000000000000; // D (0x00000000000000040000000008000000) 
14'h1301 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000001000000000000000000000000000; // D (0x00000000000000080000000008000000) 
14'h2ccc : LOC =         127'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000001000000000000000000000000000; // D (0x00000000000000100000000008000000) 
14'h1021 : LOC =         127'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000001000000000000000000000000000; // D (0x00000000000000200000000008000000) 
14'h2a8c : LOC =         127'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000001000000000000000000000000000; // D (0x00000000000000400000000008000000) 
14'h1ca1 : LOC =         127'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000001000000000000000000000000000; // D (0x00000000000000800000000008000000) 
14'h338c : LOC =         127'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000001000000000000000000000000000; // D (0x00000000000001000000000008000000) 
14'h2ea1 : LOC =         127'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000001000000000000000000000000000; // D (0x00000000000002000000000008000000) 
14'h14fb : LOC =         127'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000001000000000000000000000000000; // D (0x00000000000004000000000008000000) 
14'h2338 : LOC =         127'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000001000000000000000000000000000; // D (0x00000000000008000000000008000000) 
14'h0fc9 : LOC =         127'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000001000000000000000000000000000; // D (0x00000000000010000000000008000000) 
14'h155c : LOC =         127'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000001000000000000000000000000000; // D (0x00000000000020000000000008000000) 
14'h2076 : LOC =         127'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000001000000000000000000000000000; // D (0x00000000000040000000000008000000) 
14'h0955 : LOC =         127'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000001000000000000000000000000000; // D (0x00000000000080000000000008000000) 
14'h1864 : LOC =         127'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000001000000000000000000000000000; // D (0x00000000000100000000000008000000) 
14'h3a06 : LOC =         127'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000001000000000000000000000000000; // D (0x00000000000200000000000008000000) 
14'h3db5 : LOC =         127'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000001000000000000000000000000000; // D (0x00000000000400000000000008000000) 
14'h32d3 : LOC =         127'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000001000000000000000000000000000; // D (0x00000000000800000000000008000000) 
14'h2c1f : LOC =         127'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000001000000000000000000000000000; // D (0x00000000001000000000000008000000) 
14'h1187 : LOC =         127'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000001000000000000000000000000000; // D (0x00000000002000000000000008000000) 
14'h29c0 : LOC =         127'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000001000000000000000000000000000; // D (0x00000000004000000000000008000000) 
14'h1a39 : LOC =         127'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000001000000000000000000000000000; // D (0x00000000008000000000000008000000) 
14'h3ebc : LOC =         127'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000001000000000000000000000000000; // D (0x00000000010000000000000008000000) 
14'h34c1 : LOC =         127'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000001000000000000000000000000000; // D (0x00000000020000000000000008000000) 
14'h203b : LOC =         127'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000; // D (0x00000000040000000000000008000000) 
14'h09cf : LOC =         127'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000; // D (0x00000000080000000000000008000000) 
14'h1950 : LOC =         127'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000; // D (0x00000000100000000000000008000000) 
14'h386e : LOC =         127'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000; // D (0x00000000200000000000000008000000) 
14'h3965 : LOC =         127'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000; // D (0x00000000400000000000000008000000) 
14'h3b73 : LOC =         127'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000; // D (0x00000000800000000000000008000000) 
14'h3f5f : LOC =         127'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000; // D (0x00000001000000000000000008000000) 
14'h3707 : LOC =         127'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000; // D (0x00000002000000000000000008000000) 
14'h27b7 : LOC =         127'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000; // D (0x00000004000000000000000008000000) 
14'h06d7 : LOC =         127'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000; // D (0x00000008000000000000000008000000) 
14'h0760 : LOC =         127'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000; // D (0x00000010000000000000000008000000) 
14'h040e : LOC =         127'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000; // D (0x00000020000000000000000008000000) 
14'h02d2 : LOC =         127'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000; // D (0x00000040000000000000000008000000) 
14'h0f6a : LOC =         127'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000; // D (0x00000080000000000000000008000000) 
14'h141a : LOC =         127'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000; // D (0x00000100000000000000000008000000) 
14'h22fa : LOC =         127'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000; // D (0x00000200000000000000000008000000) 
14'h0c4d : LOC =         127'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000; // D (0x00000400000000000000000008000000) 
14'h1254 : LOC =         127'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000; // D (0x00000800000000000000000008000000) 
14'h2e66 : LOC =         127'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000; // D (0x00001000000000000000000008000000) 
14'h1575 : LOC =         127'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000; // D (0x00002000000000000000000008000000) 
14'h2024 : LOC =         127'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000; // D (0x00004000000000000000000008000000) 
14'h09f1 : LOC =         127'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000; // D (0x00008000000000000000000008000000) 
14'h192c : LOC =         127'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000; // D (0x00010000000000000000000008000000) 
14'h3896 : LOC =         127'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000; // D (0x00020000000000000000000008000000) 
14'h3895 : LOC =         127'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000; // D (0x00040000000000000000000008000000) 
14'h3893 : LOC =         127'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000; // D (0x00080000000000000000000008000000) 
14'h389f : LOC =         127'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000; // D (0x00100000000000000000000008000000) 
14'h3887 : LOC =         127'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000; // D (0x00200000000000000000000008000000) 
14'h38b7 : LOC =         127'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000; // D (0x00400000000000000000000008000000) 
14'h38d7 : LOC =         127'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000; // D (0x00800000000000000000000008000000) 
14'h3817 : LOC =         127'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000; // D (0x01000000000000000000000008000000) 
14'h3997 : LOC =         127'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000; // D (0x02000000000000000000000008000000) 
14'h3a97 : LOC =         127'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000; // D (0x04000000000000000000000008000000) 
14'h3c97 : LOC =         127'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000; // D (0x08000000000000000000000008000000) 
14'h3097 : LOC =         127'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000; // D (0x10000000000000000000000008000000) 
14'h2897 : LOC =         127'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000; // D (0x20000000000000000000000008000000) 
14'h1897 : LOC =         127'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000; // D (0x40000000000000000000000008000000) 
14'h3259 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000; // S (0x00000000000000000000000010000000) 
14'h159c : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000000000; // D (0x00000000000000000000000030000000) 
14'h3ea4 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000000000000000000000000000; // D (0x00000000000000000000000050000000) 
14'h2ba3 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000; // D (0x00000000000000000000000090000000) 
14'h01ad : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010000000000000000000000000000; // D (0x00000000000000000000000110000000) 
14'h16c6 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000010000000000000000000000000000; // D (0x00000000000000000000000210000000) 
14'h3810 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000010000000000000000000000000000; // D (0x00000000000000000000000410000000) 
14'h26cb : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000010000000000000000000000000000; // D (0x00000000000000000000000810000000) 
14'h1b7d : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000010000000000000000000000000000; // D (0x00000000000000000000001010000000) 
14'h2366 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000010000000000000000000000000000; // D (0x00000000000000000000002010000000) 
14'h1027 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000010000000000000000000000000000; // D (0x00000000000000000000004010000000) 
14'h35d2 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000010000000000000000000000000000; // D (0x00000000000000000000008010000000) 
14'h3d4f : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000010000000000000000000000000000; // D (0x00000000000000000000010010000000) 
14'h2c75 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000010000000000000000000000000000; // D (0x00000000000000000000020010000000) 
14'h0e01 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000010000000000000000000000000000; // D (0x00000000000000000000040010000000) 
14'h099e : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000010000000000000000000000000000; // D (0x00000000000000000000080010000000) 
14'h06a0 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000010000000000000000000000000000; // D (0x00000000000000000000100010000000) 
14'h18dc : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000010000000000000000000000000000; // D (0x00000000000000000000200010000000) 
14'h2424 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000010000000000000000000000000000; // D (0x00000000000000000000400010000000) 
14'h1ea3 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000010000000000000000000000000000; // D (0x00000000000000000000800010000000) 
14'h28da : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000010000000000000000000000000000; // D (0x00000000000000000001000010000000) 
14'h075f : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000010000000000000000000000000000; // D (0x00000000000000000002000010000000) 
14'h1b22 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000010000000000000000000000000000; // D (0x00000000000000000004000010000000) 
14'h23d8 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000010000000000000000000000000000; // D (0x00000000000000000008000010000000) 
14'h115b : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000010000000000000000000000000000; // D (0x00000000000000000010000010000000) 
14'h372a : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000010000000000000000000000000000; // D (0x00000000000000000020000010000000) 
14'h38bf : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000010000000000000000000000000000; // D (0x00000000000000000040000010000000) 
14'h2795 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000010000000000000000000000000000; // D (0x00000000000000000080000010000000) 
14'h19c1 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000010000000000000000000000000000; // D (0x00000000000000000100000010000000) 
14'h261e : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000010000000000000000000000000000; // D (0x00000000000000000200000010000000) 
14'h1ad7 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000010000000000000000000000000000; // D (0x00000000000000000400000010000000) 
14'h2032 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000010000000000000000000000000000; // D (0x00000000000000000800000010000000) 
14'h168f : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000010000000000000000000000000000; // D (0x00000000000000001000000010000000) 
14'h3882 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000010000000000000000000000000000; // D (0x00000000000000002000000010000000) 
14'h27ef : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000; // D (0x00000000000000004000000010000000) 
14'h1935 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000010000000000000000000000000000; // D (0x00000000000000008000000010000000) 
14'h27f6 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000010000000000000000000000000000; // D (0x00000000000000010000000010000000) 
14'h1907 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000; // D (0x00000000000000020000000010000000) 
14'h2792 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000010000000000000000000000000000; // D (0x00000000000000040000000010000000) 
14'h19cf : LOC =         127'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000010000000000000000000000000000; // D (0x00000000000000080000000010000000) 
14'h2602 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000010000000000000000000000000000; // D (0x00000000000000100000000010000000) 
14'h1aef : LOC =         127'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000010000000000000000000000000000; // D (0x00000000000000200000000010000000) 
14'h2042 : LOC =         127'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000010000000000000000000000000000; // D (0x00000000000000400000000010000000) 
14'h166f : LOC =         127'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000010000000000000000000000000000; // D (0x00000000000000800000000010000000) 
14'h3942 : LOC =         127'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000010000000000000000000000000000; // D (0x00000000000001000000000010000000) 
14'h246f : LOC =         127'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000010000000000000000000000000000; // D (0x00000000000002000000000010000000) 
14'h1e35 : LOC =         127'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000010000000000000000000000000000; // D (0x00000000000004000000000010000000) 
14'h29f6 : LOC =         127'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000010000000000000000000000000000; // D (0x00000000000008000000000010000000) 
14'h0507 : LOC =         127'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000010000000000000000000000000000; // D (0x00000000000010000000000010000000) 
14'h1f92 : LOC =         127'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000010000000000000000000000000000; // D (0x00000000000020000000000010000000) 
14'h2ab8 : LOC =         127'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000010000000000000000000000000000; // D (0x00000000000040000000000010000000) 
14'h039b : LOC =         127'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000010000000000000000000000000000; // D (0x00000000000080000000000010000000) 
14'h12aa : LOC =         127'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000010000000000000000000000000000; // D (0x00000000000100000000000010000000) 
14'h30c8 : LOC =         127'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000010000000000000000000000000000; // D (0x00000000000200000000000010000000) 
14'h377b : LOC =         127'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000010000000000000000000000000000; // D (0x00000000000400000000000010000000) 
14'h381d : LOC =         127'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000010000000000000000000000000000; // D (0x00000000000800000000000010000000) 
14'h26d1 : LOC =         127'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000010000000000000000000000000000; // D (0x00000000001000000000000010000000) 
14'h1b49 : LOC =         127'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000010000000000000000000000000000; // D (0x00000000002000000000000010000000) 
14'h230e : LOC =         127'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000010000000000000000000000000000; // D (0x00000000004000000000000010000000) 
14'h10f7 : LOC =         127'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000010000000000000000000000000000; // D (0x00000000008000000000000010000000) 
14'h3472 : LOC =         127'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000010000000000000000000000000000; // D (0x00000000010000000000000010000000) 
14'h3e0f : LOC =         127'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000010000000000000000000000000000; // D (0x00000000020000000000000010000000) 
14'h2af5 : LOC =         127'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000; // D (0x00000000040000000000000010000000) 
14'h0301 : LOC =         127'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000; // D (0x00000000080000000000000010000000) 
14'h139e : LOC =         127'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000; // D (0x00000000100000000000000010000000) 
14'h32a0 : LOC =         127'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000; // D (0x00000000200000000000000010000000) 
14'h33ab : LOC =         127'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000; // D (0x00000000400000000000000010000000) 
14'h31bd : LOC =         127'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000; // D (0x00000000800000000000000010000000) 
14'h3591 : LOC =         127'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000; // D (0x00000001000000000000000010000000) 
14'h3dc9 : LOC =         127'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000; // D (0x00000002000000000000000010000000) 
14'h2d79 : LOC =         127'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000; // D (0x00000004000000000000000010000000) 
14'h0c19 : LOC =         127'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000; // D (0x00000008000000000000000010000000) 
14'h0dae : LOC =         127'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000; // D (0x00000010000000000000000010000000) 
14'h0ec0 : LOC =         127'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000; // D (0x00000020000000000000000010000000) 
14'h081c : LOC =         127'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000; // D (0x00000040000000000000000010000000) 
14'h05a4 : LOC =         127'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000; // D (0x00000080000000000000000010000000) 
14'h1ed4 : LOC =         127'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000; // D (0x00000100000000000000000010000000) 
14'h2834 : LOC =         127'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000; // D (0x00000200000000000000000010000000) 
14'h0683 : LOC =         127'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000; // D (0x00000400000000000000000010000000) 
14'h189a : LOC =         127'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000; // D (0x00000800000000000000000010000000) 
14'h24a8 : LOC =         127'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000; // D (0x00001000000000000000000010000000) 
14'h1fbb : LOC =         127'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000; // D (0x00002000000000000000000010000000) 
14'h2aea : LOC =         127'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000; // D (0x00004000000000000000000010000000) 
14'h033f : LOC =         127'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000; // D (0x00008000000000000000000010000000) 
14'h13e2 : LOC =         127'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000; // D (0x00010000000000000000000010000000) 
14'h3258 : LOC =         127'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000; // D (0x00020000000000000000000010000000) 
14'h325b : LOC =         127'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000; // D (0x00040000000000000000000010000000) 
14'h325d : LOC =         127'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000; // D (0x00080000000000000000000010000000) 
14'h3251 : LOC =         127'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000; // D (0x00100000000000000000000010000000) 
14'h3249 : LOC =         127'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000; // D (0x00200000000000000000000010000000) 
14'h3279 : LOC =         127'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000; // D (0x00400000000000000000000010000000) 
14'h3219 : LOC =         127'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000; // D (0x00800000000000000000000010000000) 
14'h32d9 : LOC =         127'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000; // D (0x01000000000000000000000010000000) 
14'h3359 : LOC =         127'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000; // D (0x02000000000000000000000010000000) 
14'h3059 : LOC =         127'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000; // D (0x04000000000000000000000010000000) 
14'h3659 : LOC =         127'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000; // D (0x08000000000000000000000010000000) 
14'h3a59 : LOC =         127'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000; // D (0x10000000000000000000000010000000) 
14'h2259 : LOC =         127'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000; // D (0x20000000000000000000000010000000) 
14'h1259 : LOC =         127'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000; // D (0x40000000000000000000000010000000) 
14'h27c5 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000; // S (0x00000000000000000000000020000000) 
14'h2b38 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000; // D (0x00000000000000000000000060000000) 
14'h3e3f : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000000; // D (0x000000000000000000000000a0000000) 
14'h1431 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000; // D (0x00000000000000000000000120000000) 
14'h035a : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000100000000000000000000000000000; // D (0x00000000000000000000000220000000) 
14'h2d8c : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000100000000000000000000000000000; // D (0x00000000000000000000000420000000) 
14'h3357 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000100000000000000000000000000000; // D (0x00000000000000000000000820000000) 
14'h0ee1 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000100000000000000000000000000000; // D (0x00000000000000000000001020000000) 
14'h36fa : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000100000000000000000000000000000; // D (0x00000000000000000000002020000000) 
14'h05bb : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000100000000000000000000000000000; // D (0x00000000000000000000004020000000) 
14'h204e : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000100000000000000000000000000000; // D (0x00000000000000000000008020000000) 
14'h28d3 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000100000000000000000000000000000; // D (0x00000000000000000000010020000000) 
14'h39e9 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000100000000000000000000000000000; // D (0x00000000000000000000020020000000) 
14'h1b9d : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000100000000000000000000000000000; // D (0x00000000000000000000040020000000) 
14'h1c02 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000100000000000000000000000000000; // D (0x00000000000000000000080020000000) 
14'h133c : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000100000000000000000000000000000; // D (0x00000000000000000000100020000000) 
14'h0d40 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000100000000000000000000000000000; // D (0x00000000000000000000200020000000) 
14'h31b8 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000100000000000000000000000000000; // D (0x00000000000000000000400020000000) 
14'h0b3f : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000100000000000000000000000000000; // D (0x00000000000000000000800020000000) 
14'h3d46 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000100000000000000000000000000000; // D (0x00000000000000000001000020000000) 
14'h12c3 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000100000000000000000000000000000; // D (0x00000000000000000002000020000000) 
14'h0ebe : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000100000000000000000000000000000; // D (0x00000000000000000004000020000000) 
14'h3644 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000100000000000000000000000000000; // D (0x00000000000000000008000020000000) 
14'h04c7 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000100000000000000000000000000000; // D (0x00000000000000000010000020000000) 
14'h22b6 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000100000000000000000000000000000; // D (0x00000000000000000020000020000000) 
14'h2d23 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000100000000000000000000000000000; // D (0x00000000000000000040000020000000) 
14'h3209 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000100000000000000000000000000000; // D (0x00000000000000000080000020000000) 
14'h0c5d : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000100000000000000000000000000000; // D (0x00000000000000000100000020000000) 
14'h3382 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000100000000000000000000000000000; // D (0x00000000000000000200000020000000) 
14'h0f4b : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000100000000000000000000000000000; // D (0x00000000000000000400000020000000) 
14'h35ae : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000100000000000000000000000000000; // D (0x00000000000000000800000020000000) 
14'h0313 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000100000000000000000000000000000; // D (0x00000000000000001000000020000000) 
14'h2d1e : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000100000000000000000000000000000; // D (0x00000000000000002000000020000000) 
14'h3273 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000100000000000000000000000000000; // D (0x00000000000000004000000020000000) 
14'h0ca9 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000100000000000000000000000000000; // D (0x00000000000000008000000020000000) 
14'h326a : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000100000000000000000000000000000; // D (0x00000000000000010000000020000000) 
14'h0c9b : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000100000000000000000000000000000; // D (0x00000000000000020000000020000000) 
14'h320e : LOC =         127'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000100000000000000000000000000000; // D (0x00000000000000040000000020000000) 
14'h0c53 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000100000000000000000000000000000; // D (0x00000000000000080000000020000000) 
14'h339e : LOC =         127'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000100000000000000000000000000000; // D (0x00000000000000100000000020000000) 
14'h0f73 : LOC =         127'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000100000000000000000000000000000; // D (0x00000000000000200000000020000000) 
14'h35de : LOC =         127'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000100000000000000000000000000000; // D (0x00000000000000400000000020000000) 
14'h03f3 : LOC =         127'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000100000000000000000000000000000; // D (0x00000000000000800000000020000000) 
14'h2cde : LOC =         127'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000100000000000000000000000000000; // D (0x00000000000001000000000020000000) 
14'h31f3 : LOC =         127'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000100000000000000000000000000000; // D (0x00000000000002000000000020000000) 
14'h0ba9 : LOC =         127'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000100000000000000000000000000000; // D (0x00000000000004000000000020000000) 
14'h3c6a : LOC =         127'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000100000000000000000000000000000; // D (0x00000000000008000000000020000000) 
14'h109b : LOC =         127'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000100000000000000000000000000000; // D (0x00000000000010000000000020000000) 
14'h0a0e : LOC =         127'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000100000000000000000000000000000; // D (0x00000000000020000000000020000000) 
14'h3f24 : LOC =         127'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000100000000000000000000000000000; // D (0x00000000000040000000000020000000) 
14'h1607 : LOC =         127'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000100000000000000000000000000000; // D (0x00000000000080000000000020000000) 
14'h0736 : LOC =         127'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000100000000000000000000000000000; // D (0x00000000000100000000000020000000) 
14'h2554 : LOC =         127'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000100000000000000000000000000000; // D (0x00000000000200000000000020000000) 
14'h22e7 : LOC =         127'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000100000000000000000000000000000; // D (0x00000000000400000000000020000000) 
14'h2d81 : LOC =         127'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000100000000000000000000000000000; // D (0x00000000000800000000000020000000) 
14'h334d : LOC =         127'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000100000000000000000000000000000; // D (0x00000000001000000000000020000000) 
14'h0ed5 : LOC =         127'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000100000000000000000000000000000; // D (0x00000000002000000000000020000000) 
14'h3692 : LOC =         127'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000100000000000000000000000000000; // D (0x00000000004000000000000020000000) 
14'h056b : LOC =         127'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000100000000000000000000000000000; // D (0x00000000008000000000000020000000) 
14'h21ee : LOC =         127'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000100000000000000000000000000000; // D (0x00000000010000000000000020000000) 
14'h2b93 : LOC =         127'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000100000000000000000000000000000; // D (0x00000000020000000000000020000000) 
14'h3f69 : LOC =         127'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000; // D (0x00000000040000000000000020000000) 
14'h169d : LOC =         127'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000; // D (0x00000000080000000000000020000000) 
14'h0602 : LOC =         127'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000; // D (0x00000000100000000000000020000000) 
14'h273c : LOC =         127'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000; // D (0x00000000200000000000000020000000) 
14'h2637 : LOC =         127'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000; // D (0x00000000400000000000000020000000) 
14'h2421 : LOC =         127'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000; // D (0x00000000800000000000000020000000) 
14'h200d : LOC =         127'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000; // D (0x00000001000000000000000020000000) 
14'h2855 : LOC =         127'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000; // D (0x00000002000000000000000020000000) 
14'h38e5 : LOC =         127'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000; // D (0x00000004000000000000000020000000) 
14'h1985 : LOC =         127'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000; // D (0x00000008000000000000000020000000) 
14'h1832 : LOC =         127'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000; // D (0x00000010000000000000000020000000) 
14'h1b5c : LOC =         127'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000; // D (0x00000020000000000000000020000000) 
14'h1d80 : LOC =         127'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000; // D (0x00000040000000000000000020000000) 
14'h1038 : LOC =         127'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000; // D (0x00000080000000000000000020000000) 
14'h0b48 : LOC =         127'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000; // D (0x00000100000000000000000020000000) 
14'h3da8 : LOC =         127'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000; // D (0x00000200000000000000000020000000) 
14'h131f : LOC =         127'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000; // D (0x00000400000000000000000020000000) 
14'h0d06 : LOC =         127'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000; // D (0x00000800000000000000000020000000) 
14'h3134 : LOC =         127'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000; // D (0x00001000000000000000000020000000) 
14'h0a27 : LOC =         127'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000; // D (0x00002000000000000000000020000000) 
14'h3f76 : LOC =         127'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000; // D (0x00004000000000000000000020000000) 
14'h16a3 : LOC =         127'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000; // D (0x00008000000000000000000020000000) 
14'h067e : LOC =         127'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000; // D (0x00010000000000000000000020000000) 
14'h27c4 : LOC =         127'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000; // D (0x00020000000000000000000020000000) 
14'h27c7 : LOC =         127'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000; // D (0x00040000000000000000000020000000) 
14'h27c1 : LOC =         127'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000; // D (0x00080000000000000000000020000000) 
14'h27cd : LOC =         127'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000; // D (0x00100000000000000000000020000000) 
14'h27d5 : LOC =         127'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000; // D (0x00200000000000000000000020000000) 
14'h27e5 : LOC =         127'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000; // D (0x00400000000000000000000020000000) 
14'h2785 : LOC =         127'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000; // D (0x00800000000000000000000020000000) 
14'h2745 : LOC =         127'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000; // D (0x01000000000000000000000020000000) 
14'h26c5 : LOC =         127'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000; // D (0x02000000000000000000000020000000) 
14'h25c5 : LOC =         127'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000; // D (0x04000000000000000000000020000000) 
14'h23c5 : LOC =         127'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000; // D (0x08000000000000000000000020000000) 
14'h2fc5 : LOC =         127'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000; // D (0x10000000000000000000000020000000) 
14'h37c5 : LOC =         127'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000; // D (0x20000000000000000000000020000000) 
14'h07c5 : LOC =         127'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000; // D (0x40000000000000000000000020000000) 
14'h0cfd : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000; // S (0x00000000000000000000000040000000) 
14'h1507 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000000000; // D (0x000000000000000000000000c0000000) 
14'h3f09 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000000000000000000000000000000; // D (0x00000000000000000000000140000000) 
14'h2862 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000; // D (0x00000000000000000000000240000000) 
14'h06b4 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000000000000000000000000000000; // D (0x00000000000000000000000440000000) 
14'h186f : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100001000000000000000000000000000000; // D (0x00000000000000000000000840000000) 
14'h25d9 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000001000000000000000000000000000000; // D (0x00000000000000000000001040000000) 
14'h1dc2 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000001000000000000000000000000000000; // D (0x00000000000000000000002040000000) 
14'h2e83 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000001000000000000000000000000000000; // D (0x00000000000000000000004040000000) 
14'h0b76 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000001000000000000000000000000000000; // D (0x00000000000000000000008040000000) 
14'h03eb : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000001000000000000000000000000000000; // D (0x00000000000000000000010040000000) 
14'h12d1 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000001000000000000000000000000000000; // D (0x00000000000000000000020040000000) 
14'h30a5 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000001000000000000000000000000000000; // D (0x00000000000000000000040040000000) 
14'h373a : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000001000000000000000000000000000000; // D (0x00000000000000000000080040000000) 
14'h3804 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000001000000000000000000000000000000; // D (0x00000000000000000000100040000000) 
14'h2678 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000001000000000000000000000000000000; // D (0x00000000000000000000200040000000) 
14'h1a80 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001000000000000000000000000000000; // D (0x00000000000000000000400040000000) 
14'h2007 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000001000000000000000000000000000000; // D (0x00000000000000000000800040000000) 
14'h167e : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000001000000000000000000000000000000; // D (0x00000000000000000001000040000000) 
14'h39fb : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000001000000000000000000000000000000; // D (0x00000000000000000002000040000000) 
14'h2586 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000001000000000000000000000000000000; // D (0x00000000000000000004000040000000) 
14'h1d7c : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000001000000000000000000000000000000; // D (0x00000000000000000008000040000000) 
14'h2fff : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000001000000000000000000000000000000; // D (0x00000000000000000010000040000000) 
14'h098e : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000001000000000000000000000000000000; // D (0x00000000000000000020000040000000) 
14'h061b : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000001000000000000000000000000000000; // D (0x00000000000000000040000040000000) 
14'h1931 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000001000000000000000000000000000000; // D (0x00000000000000000080000040000000) 
14'h2765 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000001000000000000000000000000000000; // D (0x00000000000000000100000040000000) 
14'h18ba : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000001000000000000000000000000000000; // D (0x00000000000000000200000040000000) 
14'h2473 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000001000000000000000000000000000000; // D (0x00000000000000000400000040000000) 
14'h1e96 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000001000000000000000000000000000000; // D (0x00000000000000000800000040000000) 
14'h282b : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000001000000000000000000000000000000; // D (0x00000000000000001000000040000000) 
14'h0626 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000001000000000000000000000000000000; // D (0x00000000000000002000000040000000) 
14'h194b : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000001000000000000000000000000000000; // D (0x00000000000000004000000040000000) 
14'h2791 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000001000000000000000000000000000000; // D (0x00000000000000008000000040000000) 
14'h1952 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000; // D (0x00000000000000010000000040000000) 
14'h27a3 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000001000000000000000000000000000000; // D (0x00000000000000020000000040000000) 
14'h1936 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000001000000000000000000000000000000; // D (0x00000000000000040000000040000000) 
14'h276b : LOC =         127'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000001000000000000000000000000000000; // D (0x00000000000000080000000040000000) 
14'h18a6 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000000000000000000000000; // D (0x00000000000000100000000040000000) 
14'h244b : LOC =         127'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000001000000000000000000000000000000; // D (0x00000000000000200000000040000000) 
14'h1ee6 : LOC =         127'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000001000000000000000000000000000000; // D (0x00000000000000400000000040000000) 
14'h28cb : LOC =         127'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000001000000000000000000000000000000; // D (0x00000000000000800000000040000000) 
14'h07e6 : LOC =         127'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000001000000000000000000000000000000; // D (0x00000000000001000000000040000000) 
14'h1acb : LOC =         127'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000001000000000000000000000000000000; // D (0x00000000000002000000000040000000) 
14'h2091 : LOC =         127'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000001000000000000000000000000000000; // D (0x00000000000004000000000040000000) 
14'h1752 : LOC =         127'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000001000000000000000000000000000000; // D (0x00000000000008000000000040000000) 
14'h3ba3 : LOC =         127'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000001000000000000000000000000000000; // D (0x00000000000010000000000040000000) 
14'h2136 : LOC =         127'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000001000000000000000000000000000000; // D (0x00000000000020000000000040000000) 
14'h141c : LOC =         127'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000001000000000000000000000000000000; // D (0x00000000000040000000000040000000) 
14'h3d3f : LOC =         127'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000001000000000000000000000000000000; // D (0x00000000000080000000000040000000) 
14'h2c0e : LOC =         127'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000001000000000000000000000000000000; // D (0x00000000000100000000000040000000) 
14'h0e6c : LOC =         127'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000001000000000000000000000000000000; // D (0x00000000000200000000000040000000) 
14'h09df : LOC =         127'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000001000000000000000000000000000000; // D (0x00000000000400000000000040000000) 
14'h06b9 : LOC =         127'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000001000000000000000000000000000000; // D (0x00000000000800000000000040000000) 
14'h1875 : LOC =         127'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000001000000000000000000000000000000; // D (0x00000000001000000000000040000000) 
14'h25ed : LOC =         127'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000001000000000000000000000000000000; // D (0x00000000002000000000000040000000) 
14'h1daa : LOC =         127'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000001000000000000000000000000000000; // D (0x00000000004000000000000040000000) 
14'h2e53 : LOC =         127'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000001000000000000000000000000000000; // D (0x00000000008000000000000040000000) 
14'h0ad6 : LOC =         127'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000001000000000000000000000000000000; // D (0x00000000010000000000000040000000) 
14'h00ab : LOC =         127'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000001000000000000000000000000000000; // D (0x00000000020000000000000040000000) 
14'h1451 : LOC =         127'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000; // D (0x00000000040000000000000040000000) 
14'h3da5 : LOC =         127'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000; // D (0x00000000080000000000000040000000) 
14'h2d3a : LOC =         127'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000; // D (0x00000000100000000000000040000000) 
14'h0c04 : LOC =         127'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000; // D (0x00000000200000000000000040000000) 
14'h0d0f : LOC =         127'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000; // D (0x00000000400000000000000040000000) 
14'h0f19 : LOC =         127'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000; // D (0x00000000800000000000000040000000) 
14'h0b35 : LOC =         127'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000; // D (0x00000001000000000000000040000000) 
14'h036d : LOC =         127'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000; // D (0x00000002000000000000000040000000) 
14'h13dd : LOC =         127'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000; // D (0x00000004000000000000000040000000) 
14'h32bd : LOC =         127'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000; // D (0x00000008000000000000000040000000) 
14'h330a : LOC =         127'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000; // D (0x00000010000000000000000040000000) 
14'h3064 : LOC =         127'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000; // D (0x00000020000000000000000040000000) 
14'h36b8 : LOC =         127'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000; // D (0x00000040000000000000000040000000) 
14'h3b00 : LOC =         127'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000; // D (0x00000080000000000000000040000000) 
14'h2070 : LOC =         127'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000; // D (0x00000100000000000000000040000000) 
14'h1690 : LOC =         127'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000; // D (0x00000200000000000000000040000000) 
14'h3827 : LOC =         127'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000; // D (0x00000400000000000000000040000000) 
14'h263e : LOC =         127'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000; // D (0x00000800000000000000000040000000) 
14'h1a0c : LOC =         127'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000; // D (0x00001000000000000000000040000000) 
14'h211f : LOC =         127'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000; // D (0x00002000000000000000000040000000) 
14'h144e : LOC =         127'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000; // D (0x00004000000000000000000040000000) 
14'h3d9b : LOC =         127'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000; // D (0x00008000000000000000000040000000) 
14'h2d46 : LOC =         127'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000; // D (0x00010000000000000000000040000000) 
14'h0cfc : LOC =         127'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000; // D (0x00020000000000000000000040000000) 
14'h0cff : LOC =         127'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000; // D (0x00040000000000000000000040000000) 
14'h0cf9 : LOC =         127'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000; // D (0x00080000000000000000000040000000) 
14'h0cf5 : LOC =         127'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000; // D (0x00100000000000000000000040000000) 
14'h0ced : LOC =         127'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000; // D (0x00200000000000000000000040000000) 
14'h0cdd : LOC =         127'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000; // D (0x00400000000000000000000040000000) 
14'h0cbd : LOC =         127'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000; // D (0x00800000000000000000000040000000) 
14'h0c7d : LOC =         127'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000; // D (0x01000000000000000000000040000000) 
14'h0dfd : LOC =         127'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000; // D (0x02000000000000000000000040000000) 
14'h0efd : LOC =         127'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000; // D (0x04000000000000000000000040000000) 
14'h08fd : LOC =         127'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000; // D (0x08000000000000000000000040000000) 
14'h04fd : LOC =         127'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000; // D (0x10000000000000000000000040000000) 
14'h1cfd : LOC =         127'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000; // D (0x20000000000000000000000040000000) 
14'h2cfd : LOC =         127'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000; // D (0x40000000000000000000000040000000) 
14'h19fa : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000; // S (0x00000000000000000000000080000000) 
14'h2a0e : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000000000000; // D (0x00000000000000000000000180000000) 
14'h3d65 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000000000000000000000000000000; // D (0x00000000000000000000000280000000) 
14'h13b3 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000; // D (0x00000000000000000000000480000000) 
14'h0d68 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010000000000000000000000000000000; // D (0x00000000000000000000000880000000) 
14'h30de : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000010000000000000000000000000000000; // D (0x00000000000000000000001080000000) 
14'h08c5 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000010000000000000000000000000000000; // D (0x00000000000000000000002080000000) 
14'h3b84 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000010000000000000000000000000000000; // D (0x00000000000000000000004080000000) 
14'h1e71 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000010000000000000000000000000000000; // D (0x00000000000000000000008080000000) 
14'h16ec : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000010000000000000000000000000000000; // D (0x00000000000000000000010080000000) 
14'h07d6 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000010000000000000000000000000000000; // D (0x00000000000000000000020080000000) 
14'h25a2 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000010000000000000000000000000000000; // D (0x00000000000000000000040080000000) 
14'h223d : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000010000000000000000000000000000000; // D (0x00000000000000000000080080000000) 
14'h2d03 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000010000000000000000000000000000000; // D (0x00000000000000000000100080000000) 
14'h337f : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000010000000000000000000000000000000; // D (0x00000000000000000000200080000000) 
14'h0f87 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000010000000000000000000000000000000; // D (0x00000000000000000000400080000000) 
14'h3500 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000010000000000000000000000000000000; // D (0x00000000000000000000800080000000) 
14'h0379 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000010000000000000000000000000000000; // D (0x00000000000000000001000080000000) 
14'h2cfc : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000010000000000000000000000000000000; // D (0x00000000000000000002000080000000) 
14'h3081 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000010000000000000000000000000000000; // D (0x00000000000000000004000080000000) 
14'h087b : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000010000000000000000000000000000000; // D (0x00000000000000000008000080000000) 
14'h3af8 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000010000000000000000000000000000000; // D (0x00000000000000000010000080000000) 
14'h1c89 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000010000000000000000000000000000000; // D (0x00000000000000000020000080000000) 
14'h131c : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000010000000000000000000000000000000; // D (0x00000000000000000040000080000000) 
14'h0c36 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000010000000000000000000000000000000; // D (0x00000000000000000080000080000000) 
14'h3262 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000010000000000000000000000000000000; // D (0x00000000000000000100000080000000) 
14'h0dbd : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000010000000000000000000000000000000; // D (0x00000000000000000200000080000000) 
14'h3174 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000010000000000000000000000000000000; // D (0x00000000000000000400000080000000) 
14'h0b91 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000010000000000000000000000000000000; // D (0x00000000000000000800000080000000) 
14'h3d2c : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000010000000000000000000000000000000; // D (0x00000000000000001000000080000000) 
14'h1321 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000010000000000000000000000000000000; // D (0x00000000000000002000000080000000) 
14'h0c4c : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000010000000000000000000000000000000; // D (0x00000000000000004000000080000000) 
14'h3296 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000; // D (0x00000000000000008000000080000000) 
14'h0c55 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000010000000000000000000000000000000; // D (0x00000000000000010000000080000000) 
14'h32a4 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000; // D (0x00000000000000020000000080000000) 
14'h0c31 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000010000000000000000000000000000000; // D (0x00000000000000040000000080000000) 
14'h326c : LOC =         127'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000010000000000000000000000000000000; // D (0x00000000000000080000000080000000) 
14'h0da1 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000; // D (0x00000000000000100000000080000000) 
14'h314c : LOC =         127'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000010000000000000000000000000000000; // D (0x00000000000000200000000080000000) 
14'h0be1 : LOC =         127'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000010000000000000000000000000000000; // D (0x00000000000000400000000080000000) 
14'h3dcc : LOC =         127'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000010000000000000000000000000000000; // D (0x00000000000000800000000080000000) 
14'h12e1 : LOC =         127'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000010000000000000000000000000000000; // D (0x00000000000001000000000080000000) 
14'h0fcc : LOC =         127'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000010000000000000000000000000000000; // D (0x00000000000002000000000080000000) 
14'h3596 : LOC =         127'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000010000000000000000000000000000000; // D (0x00000000000004000000000080000000) 
14'h0255 : LOC =         127'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000010000000000000000000000000000000; // D (0x00000000000008000000000080000000) 
14'h2ea4 : LOC =         127'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000010000000000000000000000000000000; // D (0x00000000000010000000000080000000) 
14'h3431 : LOC =         127'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000010000000000000000000000000000000; // D (0x00000000000020000000000080000000) 
14'h011b : LOC =         127'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000010000000000000000000000000000000; // D (0x00000000000040000000000080000000) 
14'h2838 : LOC =         127'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000010000000000000000000000000000000; // D (0x00000000000080000000000080000000) 
14'h3909 : LOC =         127'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000010000000000000000000000000000000; // D (0x00000000000100000000000080000000) 
14'h1b6b : LOC =         127'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000010000000000000000000000000000000; // D (0x00000000000200000000000080000000) 
14'h1cd8 : LOC =         127'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000010000000000000000000000000000000; // D (0x00000000000400000000000080000000) 
14'h13be : LOC =         127'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000010000000000000000000000000000000; // D (0x00000000000800000000000080000000) 
14'h0d72 : LOC =         127'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000010000000000000000000000000000000; // D (0x00000000001000000000000080000000) 
14'h30ea : LOC =         127'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000010000000000000000000000000000000; // D (0x00000000002000000000000080000000) 
14'h08ad : LOC =         127'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000010000000000000000000000000000000; // D (0x00000000004000000000000080000000) 
14'h3b54 : LOC =         127'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000010000000000000000000000000000000; // D (0x00000000008000000000000080000000) 
14'h1fd1 : LOC =         127'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000010000000000000000000000000000000; // D (0x00000000010000000000000080000000) 
14'h15ac : LOC =         127'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000010000000000000000000000000000000; // D (0x00000000020000000000000080000000) 
14'h0156 : LOC =         127'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000; // D (0x00000000040000000000000080000000) 
14'h28a2 : LOC =         127'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000; // D (0x00000000080000000000000080000000) 
14'h383d : LOC =         127'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000; // D (0x00000000100000000000000080000000) 
14'h1903 : LOC =         127'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000; // D (0x00000000200000000000000080000000) 
14'h1808 : LOC =         127'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000; // D (0x00000000400000000000000080000000) 
14'h1a1e : LOC =         127'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000; // D (0x00000000800000000000000080000000) 
14'h1e32 : LOC =         127'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000; // D (0x00000001000000000000000080000000) 
14'h166a : LOC =         127'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000; // D (0x00000002000000000000000080000000) 
14'h06da : LOC =         127'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000; // D (0x00000004000000000000000080000000) 
14'h27ba : LOC =         127'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000; // D (0x00000008000000000000000080000000) 
14'h260d : LOC =         127'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000; // D (0x00000010000000000000000080000000) 
14'h2563 : LOC =         127'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000; // D (0x00000020000000000000000080000000) 
14'h23bf : LOC =         127'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000; // D (0x00000040000000000000000080000000) 
14'h2e07 : LOC =         127'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000; // D (0x00000080000000000000000080000000) 
14'h3577 : LOC =         127'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000; // D (0x00000100000000000000000080000000) 
14'h0397 : LOC =         127'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000; // D (0x00000200000000000000000080000000) 
14'h2d20 : LOC =         127'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000; // D (0x00000400000000000000000080000000) 
14'h3339 : LOC =         127'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000; // D (0x00000800000000000000000080000000) 
14'h0f0b : LOC =         127'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000; // D (0x00001000000000000000000080000000) 
14'h3418 : LOC =         127'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000; // D (0x00002000000000000000000080000000) 
14'h0149 : LOC =         127'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000; // D (0x00004000000000000000000080000000) 
14'h289c : LOC =         127'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000; // D (0x00008000000000000000000080000000) 
14'h3841 : LOC =         127'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000; // D (0x00010000000000000000000080000000) 
14'h19fb : LOC =         127'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000; // D (0x00020000000000000000000080000000) 
14'h19f8 : LOC =         127'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000; // D (0x00040000000000000000000080000000) 
14'h19fe : LOC =         127'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000; // D (0x00080000000000000000000080000000) 
14'h19f2 : LOC =         127'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000; // D (0x00100000000000000000000080000000) 
14'h19ea : LOC =         127'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000; // D (0x00200000000000000000000080000000) 
14'h19da : LOC =         127'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000; // D (0x00400000000000000000000080000000) 
14'h19ba : LOC =         127'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000; // D (0x00800000000000000000000080000000) 
14'h197a : LOC =         127'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000; // D (0x01000000000000000000000080000000) 
14'h18fa : LOC =         127'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000; // D (0x02000000000000000000000080000000) 
14'h1bfa : LOC =         127'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000; // D (0x04000000000000000000000080000000) 
14'h1dfa : LOC =         127'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000; // D (0x08000000000000000000000080000000) 
14'h11fa : LOC =         127'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000; // D (0x10000000000000000000000080000000) 
14'h09fa : LOC =         127'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000; // D (0x20000000000000000000000080000000) 
14'h39fa : LOC =         127'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000; // D (0x40000000000000000000000080000000) 
14'h33f4 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000; // S (0x00000000000000000000000100000000) 
14'h176b : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000000; // D (0x00000000000000000000000300000000) 
14'h39bd : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000000000; // D (0x00000000000000000000000500000000) 
14'h2766 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000; // D (0x00000000000000000000000900000000) 
14'h1ad0 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000100000000000000000000000000000000; // D (0x00000000000000000000001100000000) 
14'h22cb : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000100000000000000000000000000000000; // D (0x00000000000000000000002100000000) 
14'h118a : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000100000000000000000000000000000000; // D (0x00000000000000000000004100000000) 
14'h347f : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000100000000000000000000000000000000; // D (0x00000000000000000000008100000000) 
14'h3ce2 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000100000000000000000000000000000000; // D (0x00000000000000000000010100000000) 
14'h2dd8 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000100000000000000000000000000000000; // D (0x00000000000000000000020100000000) 
14'h0fac : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000100000000000000000000000000000000; // D (0x00000000000000000000040100000000) 
14'h0833 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000100000000000000000000000000000000; // D (0x00000000000000000000080100000000) 
14'h070d : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000100000000000000000000000000000000; // D (0x00000000000000000000100100000000) 
14'h1971 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000100000000000000000000000000000000; // D (0x00000000000000000000200100000000) 
14'h2589 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000100000000000000000000000000000000; // D (0x00000000000000000000400100000000) 
14'h1f0e : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000100000000000000000000000000000000; // D (0x00000000000000000000800100000000) 
14'h2977 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000100000000000000000000000000000000; // D (0x00000000000000000001000100000000) 
14'h06f2 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000100000000000000000000000000000000; // D (0x00000000000000000002000100000000) 
14'h1a8f : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000100000000000000000000000000000000; // D (0x00000000000000000004000100000000) 
14'h2275 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000100000000000000000000000000000000; // D (0x00000000000000000008000100000000) 
14'h10f6 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000100000000000000000000000000000000; // D (0x00000000000000000010000100000000) 
14'h3687 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000100000000000000000000000000000000; // D (0x00000000000000000020000100000000) 
14'h3912 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000100000000000000000000000000000000; // D (0x00000000000000000040000100000000) 
14'h2638 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000100000000000000000000000000000000; // D (0x00000000000000000080000100000000) 
14'h186c : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000100000000000000000000000000000000; // D (0x00000000000000000100000100000000) 
14'h27b3 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000100000000000000000000000000000000; // D (0x00000000000000000200000100000000) 
14'h1b7a : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000100000000000000000000000000000000; // D (0x00000000000000000400000100000000) 
14'h219f : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000100000000000000000000000000000000; // D (0x00000000000000000800000100000000) 
14'h1722 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000100000000000000000000000000000000; // D (0x00000000000000001000000100000000) 
14'h392f : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000100000000000000000000000000000000; // D (0x00000000000000002000000100000000) 
14'h2642 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000100000000000000000000000000000000; // D (0x00000000000000004000000100000000) 
14'h1898 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000100000000000000000000000000000000; // D (0x00000000000000008000000100000000) 
14'h265b : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000100000000000000000000000000000000; // D (0x00000000000000010000000100000000) 
14'h18aa : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000100000000000000000000000000000000; // D (0x00000000000000020000000100000000) 
14'h263f : LOC =         127'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000100000000000000000000000000000000; // D (0x00000000000000040000000100000000) 
14'h1862 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000100000000000000000000000000000000; // D (0x00000000000000080000000100000000) 
14'h27af : LOC =         127'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000100000000000000000000000000000000; // D (0x00000000000000100000000100000000) 
14'h1b42 : LOC =         127'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000100000000000000000000000000000000; // D (0x00000000000000200000000100000000) 
14'h21ef : LOC =         127'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000100000000000000000000000000000000; // D (0x00000000000000400000000100000000) 
14'h17c2 : LOC =         127'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000100000000000000000000000000000000; // D (0x00000000000000800000000100000000) 
14'h38ef : LOC =         127'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000100000000000000000000000000000000; // D (0x00000000000001000000000100000000) 
14'h25c2 : LOC =         127'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000100000000000000000000000000000000; // D (0x00000000000002000000000100000000) 
14'h1f98 : LOC =         127'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000100000000000000000000000000000000; // D (0x00000000000004000000000100000000) 
14'h285b : LOC =         127'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000100000000000000000000000000000000; // D (0x00000000000008000000000100000000) 
14'h04aa : LOC =         127'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000100000000000000000000000000000000; // D (0x00000000000010000000000100000000) 
14'h1e3f : LOC =         127'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000100000000000000000000000000000000; // D (0x00000000000020000000000100000000) 
14'h2b15 : LOC =         127'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000100000000000000000000000000000000; // D (0x00000000000040000000000100000000) 
14'h0236 : LOC =         127'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000100000000000000000000000000000000; // D (0x00000000000080000000000100000000) 
14'h1307 : LOC =         127'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000100000000000000000000000000000000; // D (0x00000000000100000000000100000000) 
14'h3165 : LOC =         127'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000100000000000000000000000000000000; // D (0x00000000000200000000000100000000) 
14'h36d6 : LOC =         127'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000100000000000000000000000000000000; // D (0x00000000000400000000000100000000) 
14'h39b0 : LOC =         127'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000100000000000000000000000000000000; // D (0x00000000000800000000000100000000) 
14'h277c : LOC =         127'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000100000000000000000000000000000000; // D (0x00000000001000000000000100000000) 
14'h1ae4 : LOC =         127'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000100000000000000000000000000000000; // D (0x00000000002000000000000100000000) 
14'h22a3 : LOC =         127'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000100000000000000000000000000000000; // D (0x00000000004000000000000100000000) 
14'h115a : LOC =         127'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000100000000000000000000000000000000; // D (0x00000000008000000000000100000000) 
14'h35df : LOC =         127'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000100000000000000000000000000000000; // D (0x00000000010000000000000100000000) 
14'h3fa2 : LOC =         127'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000100000000000000000000000000000000; // D (0x00000000020000000000000100000000) 
14'h2b58 : LOC =         127'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000; // D (0x00000000040000000000000100000000) 
14'h02ac : LOC =         127'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000; // D (0x00000000080000000000000100000000) 
14'h1233 : LOC =         127'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000; // D (0x00000000100000000000000100000000) 
14'h330d : LOC =         127'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000; // D (0x00000000200000000000000100000000) 
14'h3206 : LOC =         127'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000; // D (0x00000000400000000000000100000000) 
14'h3010 : LOC =         127'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000; // D (0x00000000800000000000000100000000) 
14'h343c : LOC =         127'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000; // D (0x00000001000000000000000100000000) 
14'h3c64 : LOC =         127'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000; // D (0x00000002000000000000000100000000) 
14'h2cd4 : LOC =         127'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000; // D (0x00000004000000000000000100000000) 
14'h0db4 : LOC =         127'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000; // D (0x00000008000000000000000100000000) 
14'h0c03 : LOC =         127'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000; // D (0x00000010000000000000000100000000) 
14'h0f6d : LOC =         127'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000; // D (0x00000020000000000000000100000000) 
14'h09b1 : LOC =         127'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000; // D (0x00000040000000000000000100000000) 
14'h0409 : LOC =         127'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000; // D (0x00000080000000000000000100000000) 
14'h1f79 : LOC =         127'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000; // D (0x00000100000000000000000100000000) 
14'h2999 : LOC =         127'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000; // D (0x00000200000000000000000100000000) 
14'h072e : LOC =         127'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000; // D (0x00000400000000000000000100000000) 
14'h1937 : LOC =         127'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000; // D (0x00000800000000000000000100000000) 
14'h2505 : LOC =         127'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000; // D (0x00001000000000000000000100000000) 
14'h1e16 : LOC =         127'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000; // D (0x00002000000000000000000100000000) 
14'h2b47 : LOC =         127'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000; // D (0x00004000000000000000000100000000) 
14'h0292 : LOC =         127'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000; // D (0x00008000000000000000000100000000) 
14'h124f : LOC =         127'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000; // D (0x00010000000000000000000100000000) 
14'h33f5 : LOC =         127'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000; // D (0x00020000000000000000000100000000) 
14'h33f6 : LOC =         127'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000; // D (0x00040000000000000000000100000000) 
14'h33f0 : LOC =         127'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000; // D (0x00080000000000000000000100000000) 
14'h33fc : LOC =         127'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000; // D (0x00100000000000000000000100000000) 
14'h33e4 : LOC =         127'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000; // D (0x00200000000000000000000100000000) 
14'h33d4 : LOC =         127'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000; // D (0x00400000000000000000000100000000) 
14'h33b4 : LOC =         127'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000; // D (0x00800000000000000000000100000000) 
14'h3374 : LOC =         127'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000; // D (0x01000000000000000000000100000000) 
14'h32f4 : LOC =         127'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000; // D (0x02000000000000000000000100000000) 
14'h31f4 : LOC =         127'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000; // D (0x04000000000000000000000100000000) 
14'h37f4 : LOC =         127'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000; // D (0x08000000000000000000000100000000) 
14'h3bf4 : LOC =         127'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000; // D (0x10000000000000000000000100000000) 
14'h23f4 : LOC =         127'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000; // D (0x20000000000000000000000100000000) 
14'h13f4 : LOC =         127'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000; // D (0x40000000000000000000000100000000) 
14'h249f : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000; // S (0x00000000000000000000000200000000) 
14'h2ed6 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000000000000; // D (0x00000000000000000000000600000000) 
14'h300d : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000000000000000000000000000000000; // D (0x00000000000000000000000a00000000) 
14'h0dbb : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000; // D (0x00000000000000000000001200000000) 
14'h35a0 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000000000000000000000000000000000; // D (0x00000000000000000000002200000000) 
14'h06e1 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100001000000000000000000000000000000000; // D (0x00000000000000000000004200000000) 
14'h2314 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000001000000000000000000000000000000000; // D (0x00000000000000000000008200000000) 
14'h2b89 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000001000000000000000000000000000000000; // D (0x00000000000000000000010200000000) 
14'h3ab3 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000001000000000000000000000000000000000; // D (0x00000000000000000000020200000000) 
14'h18c7 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000001000000000000000000000000000000000; // D (0x00000000000000000000040200000000) 
14'h1f58 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000001000000000000000000000000000000000; // D (0x00000000000000000000080200000000) 
14'h1066 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000001000000000000000000000000000000000; // D (0x00000000000000000000100200000000) 
14'h0e1a : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000001000000000000000000000000000000000; // D (0x00000000000000000000200200000000) 
14'h32e2 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000001000000000000000000000000000000000; // D (0x00000000000000000000400200000000) 
14'h0865 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000001000000000000000000000000000000000; // D (0x00000000000000000000800200000000) 
14'h3e1c : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000001000000000000000000000000000000000; // D (0x00000000000000000001000200000000) 
14'h1199 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001000000000000000000000000000000000; // D (0x00000000000000000002000200000000) 
14'h0de4 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000001000000000000000000000000000000000; // D (0x00000000000000000004000200000000) 
14'h351e : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000001000000000000000000000000000000000; // D (0x00000000000000000008000200000000) 
14'h079d : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000001000000000000000000000000000000000; // D (0x00000000000000000010000200000000) 
14'h21ec : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000001000000000000000000000000000000000; // D (0x00000000000000000020000200000000) 
14'h2e79 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000001000000000000000000000000000000000; // D (0x00000000000000000040000200000000) 
14'h3153 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000001000000000000000000000000000000000; // D (0x00000000000000000080000200000000) 
14'h0f07 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000001000000000000000000000000000000000; // D (0x00000000000000000100000200000000) 
14'h30d8 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000001000000000000000000000000000000000; // D (0x00000000000000000200000200000000) 
14'h0c11 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000001000000000000000000000000000000000; // D (0x00000000000000000400000200000000) 
14'h36f4 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000001000000000000000000000000000000000; // D (0x00000000000000000800000200000000) 
14'h0049 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000001000000000000000000000000000000000; // D (0x00000000000000001000000200000000) 
14'h2e44 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000001000000000000000000000000000000000; // D (0x00000000000000002000000200000000) 
14'h3129 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000001000000000000000000000000000000000; // D (0x00000000000000004000000200000000) 
14'h0ff3 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000001000000000000000000000000000000000; // D (0x00000000000000008000000200000000) 
14'h3130 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000001000000000000000000000000000000000; // D (0x00000000000000010000000200000000) 
14'h0fc1 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000001000000000000000000000000000000000; // D (0x00000000000000020000000200000000) 
14'h3154 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000001000000000000000000000000000000000; // D (0x00000000000000040000000200000000) 
14'h0f09 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000000; // D (0x00000000000000080000000200000000) 
14'h30c4 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000001000000000000000000000000000000000; // D (0x00000000000000100000000200000000) 
14'h0c29 : LOC =         127'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000001000000000000000000000000000000000; // D (0x00000000000000200000000200000000) 
14'h3684 : LOC =         127'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000001000000000000000000000000000000000; // D (0x00000000000000400000000200000000) 
14'h00a9 : LOC =         127'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000; // D (0x00000000000000800000000200000000) 
14'h2f84 : LOC =         127'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000001000000000000000000000000000000000; // D (0x00000000000001000000000200000000) 
14'h32a9 : LOC =         127'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000001000000000000000000000000000000000; // D (0x00000000000002000000000200000000) 
14'h08f3 : LOC =         127'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000001000000000000000000000000000000000; // D (0x00000000000004000000000200000000) 
14'h3f30 : LOC =         127'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000001000000000000000000000000000000000; // D (0x00000000000008000000000200000000) 
14'h13c1 : LOC =         127'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000001000000000000000000000000000000000; // D (0x00000000000010000000000200000000) 
14'h0954 : LOC =         127'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000001000000000000000000000000000000000; // D (0x00000000000020000000000200000000) 
14'h3c7e : LOC =         127'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000001000000000000000000000000000000000; // D (0x00000000000040000000000200000000) 
14'h155d : LOC =         127'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000001000000000000000000000000000000000; // D (0x00000000000080000000000200000000) 
14'h046c : LOC =         127'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000001000000000000000000000000000000000; // D (0x00000000000100000000000200000000) 
14'h260e : LOC =         127'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000001000000000000000000000000000000000; // D (0x00000000000200000000000200000000) 
14'h21bd : LOC =         127'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000001000000000000000000000000000000000; // D (0x00000000000400000000000200000000) 
14'h2edb : LOC =         127'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000001000000000000000000000000000000000; // D (0x00000000000800000000000200000000) 
14'h3017 : LOC =         127'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000001000000000000000000000000000000000; // D (0x00000000001000000000000200000000) 
14'h0d8f : LOC =         127'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000001000000000000000000000000000000000; // D (0x00000000002000000000000200000000) 
14'h35c8 : LOC =         127'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000001000000000000000000000000000000000; // D (0x00000000004000000000000200000000) 
14'h0631 : LOC =         127'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000001000000000000000000000000000000000; // D (0x00000000008000000000000200000000) 
14'h22b4 : LOC =         127'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000001000000000000000000000000000000000; // D (0x00000000010000000000000200000000) 
14'h28c9 : LOC =         127'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000001000000000000000000000000000000000; // D (0x00000000020000000000000200000000) 
14'h3c33 : LOC =         127'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000; // D (0x00000000040000000000000200000000) 
14'h15c7 : LOC =         127'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000; // D (0x00000000080000000000000200000000) 
14'h0558 : LOC =         127'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000; // D (0x00000000100000000000000200000000) 
14'h2466 : LOC =         127'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000; // D (0x00000000200000000000000200000000) 
14'h256d : LOC =         127'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000; // D (0x00000000400000000000000200000000) 
14'h277b : LOC =         127'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000; // D (0x00000000800000000000000200000000) 
14'h2357 : LOC =         127'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000; // D (0x00000001000000000000000200000000) 
14'h2b0f : LOC =         127'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000; // D (0x00000002000000000000000200000000) 
14'h3bbf : LOC =         127'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000; // D (0x00000004000000000000000200000000) 
14'h1adf : LOC =         127'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000; // D (0x00000008000000000000000200000000) 
14'h1b68 : LOC =         127'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000; // D (0x00000010000000000000000200000000) 
14'h1806 : LOC =         127'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000; // D (0x00000020000000000000000200000000) 
14'h1eda : LOC =         127'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000; // D (0x00000040000000000000000200000000) 
14'h1362 : LOC =         127'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000; // D (0x00000080000000000000000200000000) 
14'h0812 : LOC =         127'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000; // D (0x00000100000000000000000200000000) 
14'h3ef2 : LOC =         127'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000; // D (0x00000200000000000000000200000000) 
14'h1045 : LOC =         127'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000; // D (0x00000400000000000000000200000000) 
14'h0e5c : LOC =         127'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000; // D (0x00000800000000000000000200000000) 
14'h326e : LOC =         127'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000; // D (0x00001000000000000000000200000000) 
14'h097d : LOC =         127'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000; // D (0x00002000000000000000000200000000) 
14'h3c2c : LOC =         127'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000; // D (0x00004000000000000000000200000000) 
14'h15f9 : LOC =         127'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000; // D (0x00008000000000000000000200000000) 
14'h0524 : LOC =         127'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000; // D (0x00010000000000000000000200000000) 
14'h249e : LOC =         127'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000; // D (0x00020000000000000000000200000000) 
14'h249d : LOC =         127'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000; // D (0x00040000000000000000000200000000) 
14'h249b : LOC =         127'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000; // D (0x00080000000000000000000200000000) 
14'h2497 : LOC =         127'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000; // D (0x00100000000000000000000200000000) 
14'h248f : LOC =         127'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000; // D (0x00200000000000000000000200000000) 
14'h24bf : LOC =         127'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000; // D (0x00400000000000000000000200000000) 
14'h24df : LOC =         127'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000; // D (0x00800000000000000000000200000000) 
14'h241f : LOC =         127'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000; // D (0x01000000000000000000000200000000) 
14'h259f : LOC =         127'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000; // D (0x02000000000000000000000200000000) 
14'h269f : LOC =         127'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000; // D (0x04000000000000000000000200000000) 
14'h209f : LOC =         127'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000; // D (0x08000000000000000000000200000000) 
14'h2c9f : LOC =         127'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000; // D (0x10000000000000000000000200000000) 
14'h349f : LOC =         127'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000; // D (0x20000000000000000000000200000000) 
14'h049f : LOC =         127'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000; // D (0x40000000000000000000000200000000) 
14'h0a49 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000; // S (0x00000000000000000000000400000000) 
14'h1edb : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000000000000000; // D (0x00000000000000000000000c00000000) 
14'h236d : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000000000000000000000000000000000; // D (0x00000000000000000000001400000000) 
14'h1b76 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000; // D (0x00000000000000000000002400000000) 
14'h2837 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010000000000000000000000000000000000; // D (0x00000000000000000000004400000000) 
14'h0dc2 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000010000000000000000000000000000000000; // D (0x00000000000000000000008400000000) 
14'h055f : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000010000000000000000000000000000000000; // D (0x00000000000000000000010400000000) 
14'h1465 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000010000000000000000000000000000000000; // D (0x00000000000000000000020400000000) 
14'h3611 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000010000000000000000000000000000000000; // D (0x00000000000000000000040400000000) 
14'h318e : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000010000000000000000000000000000000000; // D (0x00000000000000000000080400000000) 
14'h3eb0 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000010000000000000000000000000000000000; // D (0x00000000000000000000100400000000) 
14'h20cc : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000010000000000000000000000000000000000; // D (0x00000000000000000000200400000000) 
14'h1c34 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000010000000000000000000000000000000000; // D (0x00000000000000000000400400000000) 
14'h26b3 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000010000000000000000000000000000000000; // D (0x00000000000000000000800400000000) 
14'h10ca : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000010000000000000000000000000000000000; // D (0x00000000000000000001000400000000) 
14'h3f4f : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000010000000000000000000000000000000000; // D (0x00000000000000000002000400000000) 
14'h2332 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000010000000000000000000000000000000000; // D (0x00000000000000000004000400000000) 
14'h1bc8 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000010000000000000000000000000000000000; // D (0x00000000000000000008000400000000) 
14'h294b : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000010000000000000000000000000000000000; // D (0x00000000000000000010000400000000) 
14'h0f3a : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000010000000000000000000000000000000000; // D (0x00000000000000000020000400000000) 
14'h00af : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000010000000000000000000000000000000000; // D (0x00000000000000000040000400000000) 
14'h1f85 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000010000000000000000000000000000000000; // D (0x00000000000000000080000400000000) 
14'h21d1 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000; // D (0x00000000000000000100000400000000) 
14'h1e0e : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000010000000000000000000000000000000000; // D (0x00000000000000000200000400000000) 
14'h22c7 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000010000000000000000000000000000000000; // D (0x00000000000000000400000400000000) 
14'h1822 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000010000000000000000000000000000000000; // D (0x00000000000000000800000400000000) 
14'h2e9f : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000010000000000000000000000000000000000; // D (0x00000000000000001000000400000000) 
14'h0092 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000010000000000000000000000000000000000; // D (0x00000000000000002000000400000000) 
14'h1fff : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000010000000000000000000000000000000000; // D (0x00000000000000004000000400000000) 
14'h2125 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000010000000000000000000000000000000000; // D (0x00000000000000008000000400000000) 
14'h1fe6 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000010000000000000000000000000000000000; // D (0x00000000000000010000000400000000) 
14'h2117 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000010000000000000000000000000000000000; // D (0x00000000000000020000000400000000) 
14'h1f82 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000000; // D (0x00000000000000040000000400000000) 
14'h21df : LOC =         127'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000010000000000000000000000000000000000; // D (0x00000000000000080000000400000000) 
14'h1e12 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000; // D (0x00000000000000100000000400000000) 
14'h22ff : LOC =         127'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000010000000000000000000000000000000000; // D (0x00000000000000200000000400000000) 
14'h1852 : LOC =         127'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000010000000000000000000000000000000000; // D (0x00000000000000400000000400000000) 
14'h2e7f : LOC =         127'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000; // D (0x00000000000000800000000400000000) 
14'h0152 : LOC =         127'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000010000000000000000000000000000000000; // D (0x00000000000001000000000400000000) 
14'h1c7f : LOC =         127'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000010000000000000000000000000000000000; // D (0x00000000000002000000000400000000) 
14'h2625 : LOC =         127'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000010000000000000000000000000000000000; // D (0x00000000000004000000000400000000) 
14'h11e6 : LOC =         127'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000010000000000000000000000000000000000; // D (0x00000000000008000000000400000000) 
14'h3d17 : LOC =         127'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000010000000000000000000000000000000000; // D (0x00000000000010000000000400000000) 
14'h2782 : LOC =         127'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000010000000000000000000000000000000000; // D (0x00000000000020000000000400000000) 
14'h12a8 : LOC =         127'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000010000000000000000000000000000000000; // D (0x00000000000040000000000400000000) 
14'h3b8b : LOC =         127'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000010000000000000000000000000000000000; // D (0x00000000000080000000000400000000) 
14'h2aba : LOC =         127'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000010000000000000000000000000000000000; // D (0x00000000000100000000000400000000) 
14'h08d8 : LOC =         127'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000010000000000000000000000000000000000; // D (0x00000000000200000000000400000000) 
14'h0f6b : LOC =         127'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000010000000000000000000000000000000000; // D (0x00000000000400000000000400000000) 
14'h000d : LOC =         127'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000010000000000000000000000000000000000; // D (0x00000000000800000000000400000000) 
14'h1ec1 : LOC =         127'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000010000000000000000000000000000000000; // D (0x00000000001000000000000400000000) 
14'h2359 : LOC =         127'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000010000000000000000000000000000000000; // D (0x00000000002000000000000400000000) 
14'h1b1e : LOC =         127'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000010000000000000000000000000000000000; // D (0x00000000004000000000000400000000) 
14'h28e7 : LOC =         127'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000010000000000000000000000000000000000; // D (0x00000000008000000000000400000000) 
14'h0c62 : LOC =         127'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000010000000000000000000000000000000000; // D (0x00000000010000000000000400000000) 
14'h061f : LOC =         127'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000010000000000000000000000000000000000; // D (0x00000000020000000000000400000000) 
14'h12e5 : LOC =         127'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000; // D (0x00000000040000000000000400000000) 
14'h3b11 : LOC =         127'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000; // D (0x00000000080000000000000400000000) 
14'h2b8e : LOC =         127'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000; // D (0x00000000100000000000000400000000) 
14'h0ab0 : LOC =         127'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000; // D (0x00000000200000000000000400000000) 
14'h0bbb : LOC =         127'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000; // D (0x00000000400000000000000400000000) 
14'h09ad : LOC =         127'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000; // D (0x00000000800000000000000400000000) 
14'h0d81 : LOC =         127'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000; // D (0x00000001000000000000000400000000) 
14'h05d9 : LOC =         127'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000; // D (0x00000002000000000000000400000000) 
14'h1569 : LOC =         127'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000; // D (0x00000004000000000000000400000000) 
14'h3409 : LOC =         127'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000; // D (0x00000008000000000000000400000000) 
14'h35be : LOC =         127'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000; // D (0x00000010000000000000000400000000) 
14'h36d0 : LOC =         127'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000; // D (0x00000020000000000000000400000000) 
14'h300c : LOC =         127'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000; // D (0x00000040000000000000000400000000) 
14'h3db4 : LOC =         127'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000; // D (0x00000080000000000000000400000000) 
14'h26c4 : LOC =         127'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000; // D (0x00000100000000000000000400000000) 
14'h1024 : LOC =         127'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000; // D (0x00000200000000000000000400000000) 
14'h3e93 : LOC =         127'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000; // D (0x00000400000000000000000400000000) 
14'h208a : LOC =         127'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000; // D (0x00000800000000000000000400000000) 
14'h1cb8 : LOC =         127'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000; // D (0x00001000000000000000000400000000) 
14'h27ab : LOC =         127'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000; // D (0x00002000000000000000000400000000) 
14'h12fa : LOC =         127'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000; // D (0x00004000000000000000000400000000) 
14'h3b2f : LOC =         127'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000; // D (0x00008000000000000000000400000000) 
14'h2bf2 : LOC =         127'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000; // D (0x00010000000000000000000400000000) 
14'h0a48 : LOC =         127'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000; // D (0x00020000000000000000000400000000) 
14'h0a4b : LOC =         127'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000; // D (0x00040000000000000000000400000000) 
14'h0a4d : LOC =         127'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000; // D (0x00080000000000000000000400000000) 
14'h0a41 : LOC =         127'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000; // D (0x00100000000000000000000400000000) 
14'h0a59 : LOC =         127'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000; // D (0x00200000000000000000000400000000) 
14'h0a69 : LOC =         127'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000; // D (0x00400000000000000000000400000000) 
14'h0a09 : LOC =         127'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000; // D (0x00800000000000000000000400000000) 
14'h0ac9 : LOC =         127'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000; // D (0x01000000000000000000000400000000) 
14'h0b49 : LOC =         127'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000; // D (0x02000000000000000000000400000000) 
14'h0849 : LOC =         127'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000; // D (0x04000000000000000000000400000000) 
14'h0e49 : LOC =         127'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000; // D (0x08000000000000000000000400000000) 
14'h0249 : LOC =         127'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000; // D (0x10000000000000000000000400000000) 
14'h1a49 : LOC =         127'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000; // D (0x20000000000000000000000400000000) 
14'h2a49 : LOC =         127'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000; // D (0x40000000000000000000000400000000) 
14'h1492 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000; // S (0x00000000000000000000000800000000) 
14'h3db6 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000000000; // D (0x00000000000000000000001800000000) 
14'h05ad : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000000000000; // D (0x00000000000000000000002800000000) 
14'h36ec : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000; // D (0x00000000000000000000004800000000) 
14'h1319 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000100000000000000000000000000000000000; // D (0x00000000000000000000008800000000) 
14'h1b84 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000100000000000000000000000000000000000; // D (0x00000000000000000000010800000000) 
14'h0abe : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000100000000000000000000000000000000000; // D (0x00000000000000000000020800000000) 
14'h28ca : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000100000000000000000000000000000000000; // D (0x00000000000000000000040800000000) 
14'h2f55 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000100000000000000000000000000000000000; // D (0x00000000000000000000080800000000) 
14'h206b : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000100000000000000000000000000000000000; // D (0x00000000000000000000100800000000) 
14'h3e17 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000100000000000000000000000000000000000; // D (0x00000000000000000000200800000000) 
14'h02ef : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000100000000000000000000000000000000000; // D (0x00000000000000000000400800000000) 
14'h3868 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000100000000000000000000000000000000000; // D (0x00000000000000000000800800000000) 
14'h0e11 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000100000000000000000000000000000000000; // D (0x00000000000000000001000800000000) 
14'h2194 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000100000000000000000000000000000000000; // D (0x00000000000000000002000800000000) 
14'h3de9 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000100000000000000000000000000000000000; // D (0x00000000000000000004000800000000) 
14'h0513 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000100000000000000000000000000000000000; // D (0x00000000000000000008000800000000) 
14'h3790 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000100000000000000000000000000000000000; // D (0x00000000000000000010000800000000) 
14'h11e1 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000100000000000000000000000000000000000; // D (0x00000000000000000020000800000000) 
14'h1e74 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000100000000000000000000000000000000000; // D (0x00000000000000000040000800000000) 
14'h015e : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000100000000000000000000000000000000000; // D (0x00000000000000000080000800000000) 
14'h3f0a : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000100000000000000000000000000000000000; // D (0x00000000000000000100000800000000) 
14'h00d5 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000100000000000000000000000000000000000; // D (0x00000000000000000200000800000000) 
14'h3c1c : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000100000000000000000000000000000000000; // D (0x00000000000000000400000800000000) 
14'h06f9 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000100000000000000000000000000000000000; // D (0x00000000000000000800000800000000) 
14'h3044 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000100000000000000000000000000000000000; // D (0x00000000000000001000000800000000) 
14'h1e49 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000100000000000000000000000000000000000; // D (0x00000000000000002000000800000000) 
14'h0124 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000100000000000000000000000000000000000; // D (0x00000000000000004000000800000000) 
14'h3ffe : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000100000000000000000000000000000000000; // D (0x00000000000000008000000800000000) 
14'h013d : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000100000000000000000000000000000000000; // D (0x00000000000000010000000800000000) 
14'h3fcc : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000100000000000000000000000000000000000; // D (0x00000000000000020000000800000000) 
14'h0159 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000100000000000000000000000000000000000; // D (0x00000000000000040000000800000000) 
14'h3f04 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000100000000000000000000000000000000000; // D (0x00000000000000080000000800000000) 
14'h00c9 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000100000000000000000000000000000000000; // D (0x00000000000000100000000800000000) 
14'h3c24 : LOC =         127'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000100000000000000000000000000000000000; // D (0x00000000000000200000000800000000) 
14'h0689 : LOC =         127'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000100000000000000000000000000000000000; // D (0x00000000000000400000000800000000) 
14'h30a4 : LOC =         127'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000100000000000000000000000000000000000; // D (0x00000000000000800000000800000000) 
14'h1f89 : LOC =         127'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000100000000000000000000000000000000000; // D (0x00000000000001000000000800000000) 
14'h02a4 : LOC =         127'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000100000000000000000000000000000000000; // D (0x00000000000002000000000800000000) 
14'h38fe : LOC =         127'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000100000000000000000000000000000000000; // D (0x00000000000004000000000800000000) 
14'h0f3d : LOC =         127'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000100000000000000000000000000000000000; // D (0x00000000000008000000000800000000) 
14'h23cc : LOC =         127'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000100000000000000000000000000000000000; // D (0x00000000000010000000000800000000) 
14'h3959 : LOC =         127'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000100000000000000000000000000000000000; // D (0x00000000000020000000000800000000) 
14'h0c73 : LOC =         127'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000100000000000000000000000000000000000; // D (0x00000000000040000000000800000000) 
14'h2550 : LOC =         127'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000100000000000000000000000000000000000; // D (0x00000000000080000000000800000000) 
14'h3461 : LOC =         127'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000100000000000000000000000000000000000; // D (0x00000000000100000000000800000000) 
14'h1603 : LOC =         127'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000100000000000000000000000000000000000; // D (0x00000000000200000000000800000000) 
14'h11b0 : LOC =         127'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000100000000000000000000000000000000000; // D (0x00000000000400000000000800000000) 
14'h1ed6 : LOC =         127'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000100000000000000000000000000000000000; // D (0x00000000000800000000000800000000) 
14'h001a : LOC =         127'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000100000000000000000000000000000000000; // D (0x00000000001000000000000800000000) 
14'h3d82 : LOC =         127'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000100000000000000000000000000000000000; // D (0x00000000002000000000000800000000) 
14'h05c5 : LOC =         127'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000100000000000000000000000000000000000; // D (0x00000000004000000000000800000000) 
14'h363c : LOC =         127'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000100000000000000000000000000000000000; // D (0x00000000008000000000000800000000) 
14'h12b9 : LOC =         127'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000100000000000000000000000000000000000; // D (0x00000000010000000000000800000000) 
14'h18c4 : LOC =         127'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000100000000000000000000000000000000000; // D (0x00000000020000000000000800000000) 
14'h0c3e : LOC =         127'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000; // D (0x00000000040000000000000800000000) 
14'h25ca : LOC =         127'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000; // D (0x00000000080000000000000800000000) 
14'h3555 : LOC =         127'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000; // D (0x00000000100000000000000800000000) 
14'h146b : LOC =         127'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000; // D (0x00000000200000000000000800000000) 
14'h1560 : LOC =         127'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000; // D (0x00000000400000000000000800000000) 
14'h1776 : LOC =         127'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000; // D (0x00000000800000000000000800000000) 
14'h135a : LOC =         127'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000; // D (0x00000001000000000000000800000000) 
14'h1b02 : LOC =         127'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000; // D (0x00000002000000000000000800000000) 
14'h0bb2 : LOC =         127'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000; // D (0x00000004000000000000000800000000) 
14'h2ad2 : LOC =         127'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000; // D (0x00000008000000000000000800000000) 
14'h2b65 : LOC =         127'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000; // D (0x00000010000000000000000800000000) 
14'h280b : LOC =         127'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000; // D (0x00000020000000000000000800000000) 
14'h2ed7 : LOC =         127'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000; // D (0x00000040000000000000000800000000) 
14'h236f : LOC =         127'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000; // D (0x00000080000000000000000800000000) 
14'h381f : LOC =         127'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000; // D (0x00000100000000000000000800000000) 
14'h0eff : LOC =         127'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000; // D (0x00000200000000000000000800000000) 
14'h2048 : LOC =         127'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000; // D (0x00000400000000000000000800000000) 
14'h3e51 : LOC =         127'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000; // D (0x00000800000000000000000800000000) 
14'h0263 : LOC =         127'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000; // D (0x00001000000000000000000800000000) 
14'h3970 : LOC =         127'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000; // D (0x00002000000000000000000800000000) 
14'h0c21 : LOC =         127'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000; // D (0x00004000000000000000000800000000) 
14'h25f4 : LOC =         127'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000; // D (0x00008000000000000000000800000000) 
14'h3529 : LOC =         127'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000; // D (0x00010000000000000000000800000000) 
14'h1493 : LOC =         127'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000; // D (0x00020000000000000000000800000000) 
14'h1490 : LOC =         127'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000; // D (0x00040000000000000000000800000000) 
14'h1496 : LOC =         127'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000; // D (0x00080000000000000000000800000000) 
14'h149a : LOC =         127'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000; // D (0x00100000000000000000000800000000) 
14'h1482 : LOC =         127'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000; // D (0x00200000000000000000000800000000) 
14'h14b2 : LOC =         127'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000; // D (0x00400000000000000000000800000000) 
14'h14d2 : LOC =         127'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000; // D (0x00800000000000000000000800000000) 
14'h1412 : LOC =         127'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000; // D (0x01000000000000000000000800000000) 
14'h1592 : LOC =         127'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000; // D (0x02000000000000000000000800000000) 
14'h1692 : LOC =         127'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000; // D (0x04000000000000000000000800000000) 
14'h1092 : LOC =         127'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000; // D (0x08000000000000000000000800000000) 
14'h1c92 : LOC =         127'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000; // D (0x10000000000000000000000800000000) 
14'h0492 : LOC =         127'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000; // D (0x20000000000000000000000800000000) 
14'h3492 : LOC =         127'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000; // D (0x40000000000000000000000800000000) 
14'h2924 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000; // S (0x00000000000000000000001000000000) 
14'h381b : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000000000000000; // D (0x00000000000000000000003000000000) 
14'h0b5a : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000000000000000000000000000000000000; // D (0x00000000000000000000005000000000) 
14'h2eaf : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000; // D (0x00000000000000000000009000000000) 
14'h2632 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000000000000000000000000000000000000; // D (0x00000000000000000000011000000000) 
14'h3708 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000100001000000000000000000000000000000000000; // D (0x00000000000000000000021000000000) 
14'h157c : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001000001000000000000000000000000000000000000; // D (0x00000000000000000000041000000000) 
14'h12e3 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010000001000000000000000000000000000000000000; // D (0x00000000000000000000081000000000) 
14'h1ddd : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100000001000000000000000000000000000000000000; // D (0x00000000000000000000101000000000) 
14'h03a1 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000000001000000000000000000000000000000000000; // D (0x00000000000000000000201000000000) 
14'h3f59 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000000001000000000000000000000000000000000000; // D (0x00000000000000000000401000000000) 
14'h05de : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000000001000000000000000000000000000000000000; // D (0x00000000000000000000801000000000) 
14'h33a7 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000000001000000000000000000000000000000000000; // D (0x00000000000000000001001000000000) 
14'h1c22 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000000001000000000000000000000000000000000000; // D (0x00000000000000000002001000000000) 
14'h005f : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000000001000000000000000000000000000000000000; // D (0x00000000000000000004001000000000) 
14'h38a5 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000000001000000000000000000000000000000000000; // D (0x00000000000000000008001000000000) 
14'h0a26 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001000000000000000000000000000000000000; // D (0x00000000000000000010001000000000) 
14'h2c57 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000000001000000000000000000000000000000000000; // D (0x00000000000000000020001000000000) 
14'h23c2 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000000001000000000000000000000000000000000000; // D (0x00000000000000000040001000000000) 
14'h3ce8 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000000001000000000000000000000000000000000000; // D (0x00000000000000000080001000000000) 
14'h02bc : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000000001000000000000000000000000000000000000; // D (0x00000000000000000100001000000000) 
14'h3d63 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000000001000000000000000000000000000000000000; // D (0x00000000000000000200001000000000) 
14'h01aa : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000000001000000000000000000000000000000000000; // D (0x00000000000000000400001000000000) 
14'h3b4f : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000000001000000000000000000000000000000000000; // D (0x00000000000000000800001000000000) 
14'h0df2 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000000001000000000000000000000000000000000000; // D (0x00000000000000001000001000000000) 
14'h23ff : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000000001000000000000000000000000000000000000; // D (0x00000000000000002000001000000000) 
14'h3c92 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000000001000000000000000000000000000000000000; // D (0x00000000000000004000001000000000) 
14'h0248 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000000001000000000000000000000000000000000000; // D (0x00000000000000008000001000000000) 
14'h3c8b : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000000001000000000000000000000000000000000000; // D (0x00000000000000010000001000000000) 
14'h027a : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000000001000000000000000000000000000000000000; // D (0x00000000000000020000001000000000) 
14'h3cef : LOC =         127'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000000001000000000000000000000000000000000000; // D (0x00000000000000040000001000000000) 
14'h02b2 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000000001000000000000000000000000000000000000; // D (0x00000000000000080000001000000000) 
14'h3d7f : LOC =         127'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000000001000000000000000000000000000000000000; // D (0x00000000000000100000001000000000) 
14'h0192 : LOC =         127'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000000001000000000000000000000000000000000000; // D (0x00000000000000200000001000000000) 
14'h3b3f : LOC =         127'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000000000; // D (0x00000000000000400000001000000000) 
14'h0d12 : LOC =         127'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000000001000000000000000000000000000000000000; // D (0x00000000000000800000001000000000) 
14'h223f : LOC =         127'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000000001000000000000000000000000000000000000; // D (0x00000000000001000000001000000000) 
14'h3f12 : LOC =         127'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000000001000000000000000000000000000000000000; // D (0x00000000000002000000001000000000) 
14'h0548 : LOC =         127'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000; // D (0x00000000000004000000001000000000) 
14'h328b : LOC =         127'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000000001000000000000000000000000000000000000; // D (0x00000000000008000000001000000000) 
14'h1e7a : LOC =         127'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000000001000000000000000000000000000000000000; // D (0x00000000000010000000001000000000) 
14'h04ef : LOC =         127'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000000001000000000000000000000000000000000000; // D (0x00000000000020000000001000000000) 
14'h31c5 : LOC =         127'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000000001000000000000000000000000000000000000; // D (0x00000000000040000000001000000000) 
14'h18e6 : LOC =         127'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000000001000000000000000000000000000000000000; // D (0x00000000000080000000001000000000) 
14'h09d7 : LOC =         127'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000000001000000000000000000000000000000000000; // D (0x00000000000100000000001000000000) 
14'h2bb5 : LOC =         127'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000000001000000000000000000000000000000000000; // D (0x00000000000200000000001000000000) 
14'h2c06 : LOC =         127'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000000001000000000000000000000000000000000000; // D (0x00000000000400000000001000000000) 
14'h2360 : LOC =         127'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000000001000000000000000000000000000000000000; // D (0x00000000000800000000001000000000) 
14'h3dac : LOC =         127'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000000001000000000000000000000000000000000000; // D (0x00000000001000000000001000000000) 
14'h0034 : LOC =         127'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000000001000000000000000000000000000000000000; // D (0x00000000002000000000001000000000) 
14'h3873 : LOC =         127'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000000001000000000000000000000000000000000000; // D (0x00000000004000000000001000000000) 
14'h0b8a : LOC =         127'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000000001000000000000000000000000000000000000; // D (0x00000000008000000000001000000000) 
14'h2f0f : LOC =         127'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000000001000000000000000000000000000000000000; // D (0x00000000010000000000001000000000) 
14'h2572 : LOC =         127'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000000001000000000000000000000000000000000000; // D (0x00000000020000000000001000000000) 
14'h3188 : LOC =         127'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000; // D (0x00000000040000000000001000000000) 
14'h187c : LOC =         127'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000; // D (0x00000000080000000000001000000000) 
14'h08e3 : LOC =         127'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000; // D (0x00000000100000000000001000000000) 
14'h29dd : LOC =         127'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000; // D (0x00000000200000000000001000000000) 
14'h28d6 : LOC =         127'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000; // D (0x00000000400000000000001000000000) 
14'h2ac0 : LOC =         127'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000; // D (0x00000000800000000000001000000000) 
14'h2eec : LOC =         127'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000; // D (0x00000001000000000000001000000000) 
14'h26b4 : LOC =         127'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000; // D (0x00000002000000000000001000000000) 
14'h3604 : LOC =         127'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000; // D (0x00000004000000000000001000000000) 
14'h1764 : LOC =         127'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000; // D (0x00000008000000000000001000000000) 
14'h16d3 : LOC =         127'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000; // D (0x00000010000000000000001000000000) 
14'h15bd : LOC =         127'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000; // D (0x00000020000000000000001000000000) 
14'h1361 : LOC =         127'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000; // D (0x00000040000000000000001000000000) 
14'h1ed9 : LOC =         127'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000; // D (0x00000080000000000000001000000000) 
14'h05a9 : LOC =         127'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000; // D (0x00000100000000000000001000000000) 
14'h3349 : LOC =         127'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000; // D (0x00000200000000000000001000000000) 
14'h1dfe : LOC =         127'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000; // D (0x00000400000000000000001000000000) 
14'h03e7 : LOC =         127'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000; // D (0x00000800000000000000001000000000) 
14'h3fd5 : LOC =         127'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000; // D (0x00001000000000000000001000000000) 
14'h04c6 : LOC =         127'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000; // D (0x00002000000000000000001000000000) 
14'h3197 : LOC =         127'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000; // D (0x00004000000000000000001000000000) 
14'h1842 : LOC =         127'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000; // D (0x00008000000000000000001000000000) 
14'h089f : LOC =         127'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000; // D (0x00010000000000000000001000000000) 
14'h2925 : LOC =         127'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000; // D (0x00020000000000000000001000000000) 
14'h2926 : LOC =         127'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000; // D (0x00040000000000000000001000000000) 
14'h2920 : LOC =         127'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000; // D (0x00080000000000000000001000000000) 
14'h292c : LOC =         127'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000; // D (0x00100000000000000000001000000000) 
14'h2934 : LOC =         127'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000; // D (0x00200000000000000000001000000000) 
14'h2904 : LOC =         127'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000; // D (0x00400000000000000000001000000000) 
14'h2964 : LOC =         127'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000; // D (0x00800000000000000000001000000000) 
14'h29a4 : LOC =         127'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000; // D (0x01000000000000000000001000000000) 
14'h2824 : LOC =         127'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000; // D (0x02000000000000000000001000000000) 
14'h2b24 : LOC =         127'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000; // D (0x04000000000000000000001000000000) 
14'h2d24 : LOC =         127'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000; // D (0x08000000000000000000001000000000) 
14'h2124 : LOC =         127'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000; // D (0x10000000000000000000001000000000) 
14'h3924 : LOC =         127'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000; // D (0x20000000000000000000001000000000) 
14'h0924 : LOC =         127'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000; // D (0x40000000000000000000001000000000) 
14'h113f : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000; // S (0x00000000000000000000002000000000) 
14'h3341 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000000000000000000; // D (0x00000000000000000000006000000000) 
14'h16b4 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000000000000000000000000000000000000; // D (0x0000000000000000000000a000000000) 
14'h1e29 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000; // D (0x00000000000000000000012000000000) 
14'h0f13 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010000000000000000000000000000000000000; // D (0x00000000000000000000022000000000) 
14'h2d67 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001000010000000000000000000000000000000000000; // D (0x00000000000000000000042000000000) 
14'h2af8 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010000010000000000000000000000000000000000000; // D (0x00000000000000000000082000000000) 
14'h25c6 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100000010000000000000000000000000000000000000; // D (0x00000000000000000000102000000000) 
14'h3bba : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000000010000000000000000000000000000000000000; // D (0x00000000000000000000202000000000) 
14'h0742 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000000010000000000000000000000000000000000000; // D (0x00000000000000000000402000000000) 
14'h3dc5 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000000010000000000000000000000000000000000000; // D (0x00000000000000000000802000000000) 
14'h0bbc : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000000010000000000000000000000000000000000000; // D (0x00000000000000000001002000000000) 
14'h2439 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000000010000000000000000000000000000000000000; // D (0x00000000000000000002002000000000) 
14'h3844 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000000010000000000000000000000000000000000000; // D (0x00000000000000000004002000000000) 
14'h00be : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000000010000000000000000000000000000000000000; // D (0x00000000000000000008002000000000) 
14'h323d : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000000010000000000000000000000000000000000000; // D (0x00000000000000000010002000000000) 
14'h144c : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000000010000000000000000000000000000000000000; // D (0x00000000000000000020002000000000) 
14'h1bd9 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000000010000000000000000000000000000000000000; // D (0x00000000000000000040002000000000) 
14'h04f3 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000000010000000000000000000000000000000000000; // D (0x00000000000000000080002000000000) 
14'h3aa7 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000000010000000000000000000000000000000000000; // D (0x00000000000000000100002000000000) 
14'h0578 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000000010000000000000000000000000000000000000; // D (0x00000000000000000200002000000000) 
14'h39b1 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000000010000000000000000000000000000000000000; // D (0x00000000000000000400002000000000) 
14'h0354 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000000; // D (0x00000000000000000800002000000000) 
14'h35e9 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000000010000000000000000000000000000000000000; // D (0x00000000000000001000002000000000) 
14'h1be4 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000000010000000000000000000000000000000000000; // D (0x00000000000000002000002000000000) 
14'h0489 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000000010000000000000000000000000000000000000; // D (0x00000000000000004000002000000000) 
14'h3a53 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000000010000000000000000000000000000000000000; // D (0x00000000000000008000002000000000) 
14'h0490 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000000010000000000000000000000000000000000000; // D (0x00000000000000010000002000000000) 
14'h3a61 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000000010000000000000000000000000000000000000; // D (0x00000000000000020000002000000000) 
14'h04f4 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000000010000000000000000000000000000000000000; // D (0x00000000000000040000002000000000) 
14'h3aa9 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000000010000000000000000000000000000000000000; // D (0x00000000000000080000002000000000) 
14'h0564 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000000010000000000000000000000000000000000000; // D (0x00000000000000100000002000000000) 
14'h3989 : LOC =         127'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000000000; // D (0x00000000000000200000002000000000) 
14'h0324 : LOC =         127'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000000010000000000000000000000000000000000000; // D (0x00000000000000400000002000000000) 
14'h3509 : LOC =         127'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000000; // D (0x00000000000000800000002000000000) 
14'h1a24 : LOC =         127'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000000010000000000000000000000000000000000000; // D (0x00000000000001000000002000000000) 
14'h0709 : LOC =         127'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000000010000000000000000000000000000000000000; // D (0x00000000000002000000002000000000) 
14'h3d53 : LOC =         127'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000000; // D (0x00000000000004000000002000000000) 
14'h0a90 : LOC =         127'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000000010000000000000000000000000000000000000; // D (0x00000000000008000000002000000000) 
14'h2661 : LOC =         127'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000000010000000000000000000000000000000000000; // D (0x00000000000010000000002000000000) 
14'h3cf4 : LOC =         127'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000000010000000000000000000000000000000000000; // D (0x00000000000020000000002000000000) 
14'h09de : LOC =         127'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000000010000000000000000000000000000000000000; // D (0x00000000000040000000002000000000) 
14'h20fd : LOC =         127'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000000010000000000000000000000000000000000000; // D (0x00000000000080000000002000000000) 
14'h31cc : LOC =         127'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000000010000000000000000000000000000000000000; // D (0x00000000000100000000002000000000) 
14'h13ae : LOC =         127'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000000010000000000000000000000000000000000000; // D (0x00000000000200000000002000000000) 
14'h141d : LOC =         127'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000000010000000000000000000000000000000000000; // D (0x00000000000400000000002000000000) 
14'h1b7b : LOC =         127'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000000010000000000000000000000000000000000000; // D (0x00000000000800000000002000000000) 
14'h05b7 : LOC =         127'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000000010000000000000000000000000000000000000; // D (0x00000000001000000000002000000000) 
14'h382f : LOC =         127'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000000010000000000000000000000000000000000000; // D (0x00000000002000000000002000000000) 
14'h0068 : LOC =         127'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000000010000000000000000000000000000000000000; // D (0x00000000004000000000002000000000) 
14'h3391 : LOC =         127'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000000010000000000000000000000000000000000000; // D (0x00000000008000000000002000000000) 
14'h1714 : LOC =         127'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000000010000000000000000000000000000000000000; // D (0x00000000010000000000002000000000) 
14'h1d69 : LOC =         127'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000000010000000000000000000000000000000000000; // D (0x00000000020000000000002000000000) 
14'h0993 : LOC =         127'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000; // D (0x00000000040000000000002000000000) 
14'h2067 : LOC =         127'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000; // D (0x00000000080000000000002000000000) 
14'h30f8 : LOC =         127'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000; // D (0x00000000100000000000002000000000) 
14'h11c6 : LOC =         127'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000; // D (0x00000000200000000000002000000000) 
14'h10cd : LOC =         127'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000; // D (0x00000000400000000000002000000000) 
14'h12db : LOC =         127'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000; // D (0x00000000800000000000002000000000) 
14'h16f7 : LOC =         127'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000; // D (0x00000001000000000000002000000000) 
14'h1eaf : LOC =         127'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000; // D (0x00000002000000000000002000000000) 
14'h0e1f : LOC =         127'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000; // D (0x00000004000000000000002000000000) 
14'h2f7f : LOC =         127'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000; // D (0x00000008000000000000002000000000) 
14'h2ec8 : LOC =         127'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000; // D (0x00000010000000000000002000000000) 
14'h2da6 : LOC =         127'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000; // D (0x00000020000000000000002000000000) 
14'h2b7a : LOC =         127'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000; // D (0x00000040000000000000002000000000) 
14'h26c2 : LOC =         127'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000; // D (0x00000080000000000000002000000000) 
14'h3db2 : LOC =         127'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000; // D (0x00000100000000000000002000000000) 
14'h0b52 : LOC =         127'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000; // D (0x00000200000000000000002000000000) 
14'h25e5 : LOC =         127'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000; // D (0x00000400000000000000002000000000) 
14'h3bfc : LOC =         127'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000; // D (0x00000800000000000000002000000000) 
14'h07ce : LOC =         127'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000; // D (0x00001000000000000000002000000000) 
14'h3cdd : LOC =         127'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000; // D (0x00002000000000000000002000000000) 
14'h098c : LOC =         127'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000; // D (0x00004000000000000000002000000000) 
14'h2059 : LOC =         127'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000; // D (0x00008000000000000000002000000000) 
14'h3084 : LOC =         127'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000; // D (0x00010000000000000000002000000000) 
14'h113e : LOC =         127'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000; // D (0x00020000000000000000002000000000) 
14'h113d : LOC =         127'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000; // D (0x00040000000000000000002000000000) 
14'h113b : LOC =         127'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000; // D (0x00080000000000000000002000000000) 
14'h1137 : LOC =         127'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000; // D (0x00100000000000000000002000000000) 
14'h112f : LOC =         127'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000; // D (0x00200000000000000000002000000000) 
14'h111f : LOC =         127'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000; // D (0x00400000000000000000002000000000) 
14'h117f : LOC =         127'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000; // D (0x00800000000000000000002000000000) 
14'h11bf : LOC =         127'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000; // D (0x01000000000000000000002000000000) 
14'h103f : LOC =         127'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000; // D (0x02000000000000000000002000000000) 
14'h133f : LOC =         127'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000; // D (0x04000000000000000000002000000000) 
14'h153f : LOC =         127'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000; // D (0x08000000000000000000002000000000) 
14'h193f : LOC =         127'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000; // D (0x10000000000000000000002000000000) 
14'h013f : LOC =         127'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000; // D (0x20000000000000000000002000000000) 
14'h313f : LOC =         127'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000; // D (0x40000000000000000000002000000000) 
14'h227e : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000; // S (0x00000000000000000000004000000000) 
14'h25f5 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000000000000; // D (0x0000000000000000000000c000000000) 
14'h2d68 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000000000000000; // D (0x00000000000000000000014000000000) 
14'h3c52 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000; // D (0x00000000000000000000024000000000) 
14'h1e26 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001000100000000000000000000000000000000000000; // D (0x00000000000000000000044000000000) 
14'h19b9 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010000100000000000000000000000000000000000000; // D (0x00000000000000000000084000000000) 
14'h1687 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100000100000000000000000000000000000000000000; // D (0x00000000000000000000104000000000) 
14'h08fb : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000000100000000000000000000000000000000000000; // D (0x00000000000000000000204000000000) 
14'h3403 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000000100000000000000000000000000000000000000; // D (0x00000000000000000000404000000000) 
14'h0e84 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000000100000000000000000000000000000000000000; // D (0x00000000000000000000804000000000) 
14'h38fd : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000000100000000000000000000000000000000000000; // D (0x00000000000000000001004000000000) 
14'h1778 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000000100000000000000000000000000000000000000; // D (0x00000000000000000002004000000000) 
14'h0b05 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000000100000000000000000000000000000000000000; // D (0x00000000000000000004004000000000) 
14'h33ff : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000000100000000000000000000000000000000000000; // D (0x00000000000000000008004000000000) 
14'h017c : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000000100000000000000000000000000000000000000; // D (0x00000000000000000010004000000000) 
14'h270d : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000000100000000000000000000000000000000000000; // D (0x00000000000000000020004000000000) 
14'h2898 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000000100000000000000000000000000000000000000; // D (0x00000000000000000040004000000000) 
14'h37b2 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000000100000000000000000000000000000000000000; // D (0x00000000000000000080004000000000) 
14'h09e6 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000000100000000000000000000000000000000000000; // D (0x00000000000000000100004000000000) 
14'h3639 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000000100000000000000000000000000000000000000; // D (0x00000000000000000200004000000000) 
14'h0af0 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000000100000000000000000000000000000000000000; // D (0x00000000000000000400004000000000) 
14'h3015 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000000100000000000000000000000000000000000000; // D (0x00000000000000000800004000000000) 
14'h06a8 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000000100000000000000000000000000000000000000; // D (0x00000000000000001000004000000000) 
14'h28a5 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000000100000000000000000000000000000000000000; // D (0x00000000000000002000004000000000) 
14'h37c8 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000000100000000000000000000000000000000000000; // D (0x00000000000000004000004000000000) 
14'h0912 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000000100000000000000000000000000000000000000; // D (0x00000000000000008000004000000000) 
14'h37d1 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000000100000000000000000000000000000000000000; // D (0x00000000000000010000004000000000) 
14'h0920 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000000100000000000000000000000000000000000000; // D (0x00000000000000020000004000000000) 
14'h37b5 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000000100000000000000000000000000000000000000; // D (0x00000000000000040000004000000000) 
14'h09e8 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000000100000000000000000000000000000000000000; // D (0x00000000000000080000004000000000) 
14'h3625 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000000100000000000000000000000000000000000000; // D (0x00000000000000100000004000000000) 
14'h0ac8 : LOC =         127'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000000100000000000000000000000000000000000000; // D (0x00000000000000200000004000000000) 
14'h3065 : LOC =         127'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000000100000000000000000000000000000000000000; // D (0x00000000000000400000004000000000) 
14'h0648 : LOC =         127'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000000100000000000000000000000000000000000000; // D (0x00000000000000800000004000000000) 
14'h2965 : LOC =         127'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000000100000000000000000000000000000000000000; // D (0x00000000000001000000004000000000) 
14'h3448 : LOC =         127'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000000100000000000000000000000000000000000000; // D (0x00000000000002000000004000000000) 
14'h0e12 : LOC =         127'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000000100000000000000000000000000000000000000; // D (0x00000000000004000000004000000000) 
14'h39d1 : LOC =         127'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000000100000000000000000000000000000000000000; // D (0x00000000000008000000004000000000) 
14'h1520 : LOC =         127'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000000100000000000000000000000000000000000000; // D (0x00000000000010000000004000000000) 
14'h0fb5 : LOC =         127'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000000100000000000000000000000000000000000000; // D (0x00000000000020000000004000000000) 
14'h3a9f : LOC =         127'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000000100000000000000000000000000000000000000; // D (0x00000000000040000000004000000000) 
14'h13bc : LOC =         127'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000000100000000000000000000000000000000000000; // D (0x00000000000080000000004000000000) 
14'h028d : LOC =         127'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000000100000000000000000000000000000000000000; // D (0x00000000000100000000004000000000) 
14'h20ef : LOC =         127'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000000100000000000000000000000000000000000000; // D (0x00000000000200000000004000000000) 
14'h275c : LOC =         127'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000000100000000000000000000000000000000000000; // D (0x00000000000400000000004000000000) 
14'h283a : LOC =         127'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000000100000000000000000000000000000000000000; // D (0x00000000000800000000004000000000) 
14'h36f6 : LOC =         127'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000000100000000000000000000000000000000000000; // D (0x00000000001000000000004000000000) 
14'h0b6e : LOC =         127'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000000100000000000000000000000000000000000000; // D (0x00000000002000000000004000000000) 
14'h3329 : LOC =         127'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000000100000000000000000000000000000000000000; // D (0x00000000004000000000004000000000) 
14'h00d0 : LOC =         127'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000000100000000000000000000000000000000000000; // D (0x00000000008000000000004000000000) 
14'h2455 : LOC =         127'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000000100000000000000000000000000000000000000; // D (0x00000000010000000000004000000000) 
14'h2e28 : LOC =         127'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000000100000000000000000000000000000000000000; // D (0x00000000020000000000004000000000) 
14'h3ad2 : LOC =         127'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000; // D (0x00000000040000000000004000000000) 
14'h1326 : LOC =         127'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000; // D (0x00000000080000000000004000000000) 
14'h03b9 : LOC =         127'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000; // D (0x00000000100000000000004000000000) 
14'h2287 : LOC =         127'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000; // D (0x00000000200000000000004000000000) 
14'h238c : LOC =         127'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000; // D (0x00000000400000000000004000000000) 
14'h219a : LOC =         127'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000; // D (0x00000000800000000000004000000000) 
14'h25b6 : LOC =         127'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000; // D (0x00000001000000000000004000000000) 
14'h2dee : LOC =         127'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000; // D (0x00000002000000000000004000000000) 
14'h3d5e : LOC =         127'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000; // D (0x00000004000000000000004000000000) 
14'h1c3e : LOC =         127'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000; // D (0x00000008000000000000004000000000) 
14'h1d89 : LOC =         127'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000; // D (0x00000010000000000000004000000000) 
14'h1ee7 : LOC =         127'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000; // D (0x00000020000000000000004000000000) 
14'h183b : LOC =         127'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000; // D (0x00000040000000000000004000000000) 
14'h1583 : LOC =         127'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000; // D (0x00000080000000000000004000000000) 
14'h0ef3 : LOC =         127'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000; // D (0x00000100000000000000004000000000) 
14'h3813 : LOC =         127'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000; // D (0x00000200000000000000004000000000) 
14'h16a4 : LOC =         127'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000; // D (0x00000400000000000000004000000000) 
14'h08bd : LOC =         127'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000; // D (0x00000800000000000000004000000000) 
14'h348f : LOC =         127'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000; // D (0x00001000000000000000004000000000) 
14'h0f9c : LOC =         127'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000; // D (0x00002000000000000000004000000000) 
14'h3acd : LOC =         127'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000; // D (0x00004000000000000000004000000000) 
14'h1318 : LOC =         127'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000; // D (0x00008000000000000000004000000000) 
14'h03c5 : LOC =         127'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000; // D (0x00010000000000000000004000000000) 
14'h227f : LOC =         127'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000; // D (0x00020000000000000000004000000000) 
14'h227c : LOC =         127'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000; // D (0x00040000000000000000004000000000) 
14'h227a : LOC =         127'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000; // D (0x00080000000000000000004000000000) 
14'h2276 : LOC =         127'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000; // D (0x00100000000000000000004000000000) 
14'h226e : LOC =         127'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000; // D (0x00200000000000000000004000000000) 
14'h225e : LOC =         127'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000; // D (0x00400000000000000000004000000000) 
14'h223e : LOC =         127'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000; // D (0x00800000000000000000004000000000) 
14'h22fe : LOC =         127'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000; // D (0x01000000000000000000004000000000) 
14'h237e : LOC =         127'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000; // D (0x02000000000000000000004000000000) 
14'h207e : LOC =         127'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000; // D (0x04000000000000000000004000000000) 
14'h267e : LOC =         127'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000; // D (0x08000000000000000000004000000000) 
14'h2a7e : LOC =         127'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000; // D (0x10000000000000000000004000000000) 
14'h327e : LOC =         127'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000; // D (0x20000000000000000000004000000000) 
14'h027e : LOC =         127'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000; // D (0x40000000000000000000004000000000) 
14'h078b : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000; // S (0x00000000000000000000008000000000) 
14'h089d : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000000000000000000; // D (0x00000000000000000000018000000000) 
14'h19a7 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000000000000000000000000000000000000000; // D (0x00000000000000000000028000000000) 
14'h3bd3 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000; // D (0x00000000000000000000048000000000) 
14'h3c4c : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000000000000000000000000000000000000000; // D (0x00000000000000000000088000000000) 
14'h3372 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100001000000000000000000000000000000000000000; // D (0x00000000000000000000108000000000) 
14'h2d0e : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000001000000000000000000000000000000000000000; // D (0x00000000000000000000208000000000) 
14'h11f6 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000001000000000000000000000000000000000000000; // D (0x00000000000000000000408000000000) 
14'h2b71 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000001000000000000000000000000000000000000000; // D (0x00000000000000000000808000000000) 
14'h1d08 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000001000000000000000000000000000000000000000; // D (0x00000000000000000001008000000000) 
14'h328d : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000001000000000000000000000000000000000000000; // D (0x00000000000000000002008000000000) 
14'h2ef0 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000001000000000000000000000000000000000000000; // D (0x00000000000000000004008000000000) 
14'h160a : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000001000000000000000000000000000000000000000; // D (0x00000000000000000008008000000000) 
14'h2489 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000001000000000000000000000000000000000000000; // D (0x00000000000000000010008000000000) 
14'h02f8 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000001000000000000000000000000000000000000000; // D (0x00000000000000000020008000000000) 
14'h0d6d : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000001000000000000000000000000000000000000000; // D (0x00000000000000000040008000000000) 
14'h1247 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000001000000000000000000000000000000000000000; // D (0x00000000000000000080008000000000) 
14'h2c13 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000001000000000000000000000000000000000000000; // D (0x00000000000000000100008000000000) 
14'h13cc : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000001000000000000000000000000000000000000000; // D (0x00000000000000000200008000000000) 
14'h2f05 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000001000000000000000000000000000000000000000; // D (0x00000000000000000400008000000000) 
14'h15e0 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000001000000000000000000000000000000000000000; // D (0x00000000000000000800008000000000) 
14'h235d : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000001000000000000000000000000000000000000000; // D (0x00000000000000001000008000000000) 
14'h0d50 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000001000000000000000000000000000000000000000; // D (0x00000000000000002000008000000000) 
14'h123d : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000001000000000000000000000000000000000000000; // D (0x00000000000000004000008000000000) 
14'h2ce7 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000001000000000000000000000000000000000000000; // D (0x00000000000000008000008000000000) 
14'h1224 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000001000000000000000000000000000000000000000; // D (0x00000000000000010000008000000000) 
14'h2cd5 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000001000000000000000000000000000000000000000; // D (0x00000000000000020000008000000000) 
14'h1240 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000001000000000000000000000000000000000000000; // D (0x00000000000000040000008000000000) 
14'h2c1d : LOC =         127'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000001000000000000000000000000000000000000000; // D (0x00000000000000080000008000000000) 
14'h13d0 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000001000000000000000000000000000000000000000; // D (0x00000000000000100000008000000000) 
14'h2f3d : LOC =         127'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000001000000000000000000000000000000000000000; // D (0x00000000000000200000008000000000) 
14'h1590 : LOC =         127'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000001000000000000000000000000000000000000000; // D (0x00000000000000400000008000000000) 
14'h23bd : LOC =         127'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000001000000000000000000000000000000000000000; // D (0x00000000000000800000008000000000) 
14'h0c90 : LOC =         127'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000001000000000000000000000000000000000000000; // D (0x00000000000001000000008000000000) 
14'h11bd : LOC =         127'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000000000000; // D (0x00000000000002000000008000000000) 
14'h2be7 : LOC =         127'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000001000000000000000000000000000000000000000; // D (0x00000000000004000000008000000000) 
14'h1c24 : LOC =         127'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000001000000000000000000000000000000000000000; // D (0x00000000000008000000008000000000) 
14'h30d5 : LOC =         127'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000001000000000000000000000000000000000000000; // D (0x00000000000010000000008000000000) 
14'h2a40 : LOC =         127'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000000; // D (0x00000000000020000000008000000000) 
14'h1f6a : LOC =         127'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000001000000000000000000000000000000000000000; // D (0x00000000000040000000008000000000) 
14'h3649 : LOC =         127'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000001000000000000000000000000000000000000000; // D (0x00000000000080000000008000000000) 
14'h2778 : LOC =         127'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000001000000000000000000000000000000000000000; // D (0x00000000000100000000008000000000) 
14'h051a : LOC =         127'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000001000000000000000000000000000000000000000; // D (0x00000000000200000000008000000000) 
14'h02a9 : LOC =         127'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000001000000000000000000000000000000000000000; // D (0x00000000000400000000008000000000) 
14'h0dcf : LOC =         127'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000001000000000000000000000000000000000000000; // D (0x00000000000800000000008000000000) 
14'h1303 : LOC =         127'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000001000000000000000000000000000000000000000; // D (0x00000000001000000000008000000000) 
14'h2e9b : LOC =         127'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000001000000000000000000000000000000000000000; // D (0x00000000002000000000008000000000) 
14'h16dc : LOC =         127'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000001000000000000000000000000000000000000000; // D (0x00000000004000000000008000000000) 
14'h2525 : LOC =         127'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000001000000000000000000000000000000000000000; // D (0x00000000008000000000008000000000) 
14'h01a0 : LOC =         127'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000001000000000000000000000000000000000000000; // D (0x00000000010000000000008000000000) 
14'h0bdd : LOC =         127'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000001000000000000000000000000000000000000000; // D (0x00000000020000000000008000000000) 
14'h1f27 : LOC =         127'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000; // D (0x00000000040000000000008000000000) 
14'h36d3 : LOC =         127'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000; // D (0x00000000080000000000008000000000) 
14'h264c : LOC =         127'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000; // D (0x00000000100000000000008000000000) 
14'h0772 : LOC =         127'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000; // D (0x00000000200000000000008000000000) 
14'h0679 : LOC =         127'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000; // D (0x00000000400000000000008000000000) 
14'h046f : LOC =         127'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000; // D (0x00000000800000000000008000000000) 
14'h0043 : LOC =         127'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000; // D (0x00000001000000000000008000000000) 
14'h081b : LOC =         127'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000; // D (0x00000002000000000000008000000000) 
14'h18ab : LOC =         127'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000; // D (0x00000004000000000000008000000000) 
14'h39cb : LOC =         127'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000; // D (0x00000008000000000000008000000000) 
14'h387c : LOC =         127'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000; // D (0x00000010000000000000008000000000) 
14'h3b12 : LOC =         127'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000; // D (0x00000020000000000000008000000000) 
14'h3dce : LOC =         127'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000; // D (0x00000040000000000000008000000000) 
14'h3076 : LOC =         127'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000; // D (0x00000080000000000000008000000000) 
14'h2b06 : LOC =         127'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000; // D (0x00000100000000000000008000000000) 
14'h1de6 : LOC =         127'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000; // D (0x00000200000000000000008000000000) 
14'h3351 : LOC =         127'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000; // D (0x00000400000000000000008000000000) 
14'h2d48 : LOC =         127'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000; // D (0x00000800000000000000008000000000) 
14'h117a : LOC =         127'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000; // D (0x00001000000000000000008000000000) 
14'h2a69 : LOC =         127'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000; // D (0x00002000000000000000008000000000) 
14'h1f38 : LOC =         127'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000; // D (0x00004000000000000000008000000000) 
14'h36ed : LOC =         127'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000; // D (0x00008000000000000000008000000000) 
14'h2630 : LOC =         127'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000; // D (0x00010000000000000000008000000000) 
14'h078a : LOC =         127'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000; // D (0x00020000000000000000008000000000) 
14'h0789 : LOC =         127'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000; // D (0x00040000000000000000008000000000) 
14'h078f : LOC =         127'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000; // D (0x00080000000000000000008000000000) 
14'h0783 : LOC =         127'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000; // D (0x00100000000000000000008000000000) 
14'h079b : LOC =         127'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000; // D (0x00200000000000000000008000000000) 
14'h07ab : LOC =         127'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000; // D (0x00400000000000000000008000000000) 
14'h07cb : LOC =         127'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000; // D (0x00800000000000000000008000000000) 
14'h070b : LOC =         127'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000; // D (0x01000000000000000000008000000000) 
14'h068b : LOC =         127'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000; // D (0x02000000000000000000008000000000) 
14'h058b : LOC =         127'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000; // D (0x04000000000000000000008000000000) 
14'h038b : LOC =         127'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000; // D (0x08000000000000000000008000000000) 
14'h0f8b : LOC =         127'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000; // D (0x10000000000000000000008000000000) 
14'h178b : LOC =         127'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000; // D (0x20000000000000000000008000000000) 
14'h278b : LOC =         127'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000; // D (0x40000000000000000000008000000000) 
14'h0f16 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000; // S (0x00000000000000000000010000000000) 
14'h113a : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000000000000000000000; // D (0x00000000000000000000030000000000) 
14'h334e : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000000000000000000000000000000000000000; // D (0x00000000000000000000050000000000) 
14'h34d1 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000; // D (0x00000000000000000000090000000000) 
14'h3bef : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100010000000000000000000000000000000000000000; // D (0x00000000000000000000110000000000) 
14'h2593 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000010000000000000000000000000000000000000000; // D (0x00000000000000000000210000000000) 
14'h196b : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000010000000000000000000000000000000000000000; // D (0x00000000000000000000410000000000) 
14'h23ec : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000010000000000000000000000000000000000000000; // D (0x00000000000000000000810000000000) 
14'h1595 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000010000000000000000000000000000000000000000; // D (0x00000000000000000001010000000000) 
14'h3a10 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000010000000000000000000000000000000000000000; // D (0x00000000000000000002010000000000) 
14'h266d : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000010000000000000000000000000000000000000000; // D (0x00000000000000000004010000000000) 
14'h1e97 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000010000000000000000000000000000000000000000; // D (0x00000000000000000008010000000000) 
14'h2c14 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000010000000000000000000000000000000000000000; // D (0x00000000000000000010010000000000) 
14'h0a65 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000010000000000000000000000000000000000000000; // D (0x00000000000000000020010000000000) 
14'h05f0 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000010000000000000000000000000000000000000000; // D (0x00000000000000000040010000000000) 
14'h1ada : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000010000000000000000000000000000000000000000; // D (0x00000000000000000080010000000000) 
14'h248e : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000010000000000000000000000000000000000000000; // D (0x00000000000000000100010000000000) 
14'h1b51 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000010000000000000000000000000000000000000000; // D (0x00000000000000000200010000000000) 
14'h2798 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000010000000000000000000000000000000000000000; // D (0x00000000000000000400010000000000) 
14'h1d7d : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000010000000000000000000000000000000000000000; // D (0x00000000000000000800010000000000) 
14'h2bc0 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000010000000000000000000000000000000000000000; // D (0x00000000000000001000010000000000) 
14'h05cd : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000010000000000000000000000000000000000000000; // D (0x00000000000000002000010000000000) 
14'h1aa0 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000000000; // D (0x00000000000000004000010000000000) 
14'h247a : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000010000000000000000000000000000000000000000; // D (0x00000000000000008000010000000000) 
14'h1ab9 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000010000000000000000000000000000000000000000; // D (0x00000000000000010000010000000000) 
14'h2448 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000010000000000000000000000000000000000000000; // D (0x00000000000000020000010000000000) 
14'h1add : LOC =         127'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000010000000000000000000000000000000000000000; // D (0x00000000000000040000010000000000) 
14'h2480 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000010000000000000000000000000000000000000000; // D (0x00000000000000080000010000000000) 
14'h1b4d : LOC =         127'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000010000000000000000000000000000000000000000; // D (0x00000000000000100000010000000000) 
14'h27a0 : LOC =         127'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000010000000000000000000000000000000000000000; // D (0x00000000000000200000010000000000) 
14'h1d0d : LOC =         127'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000010000000000000000000000000000000000000000; // D (0x00000000000000400000010000000000) 
14'h2b20 : LOC =         127'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000010000000000000000000000000000000000000000; // D (0x00000000000000800000010000000000) 
14'h040d : LOC =         127'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000000000000; // D (0x00000000000001000000010000000000) 
14'h1920 : LOC =         127'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000010000000000000000000000000000000000000000; // D (0x00000000000002000000010000000000) 
14'h237a : LOC =         127'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000000000; // D (0x00000000000004000000010000000000) 
14'h14b9 : LOC =         127'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000010000000000000000000000000000000000000000; // D (0x00000000000008000000010000000000) 
14'h3848 : LOC =         127'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000010000000000000000000000000000000000000000; // D (0x00000000000010000000010000000000) 
14'h22dd : LOC =         127'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000000000; // D (0x00000000000020000000010000000000) 
14'h17f7 : LOC =         127'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000010000000000000000000000000000000000000000; // D (0x00000000000040000000010000000000) 
14'h3ed4 : LOC =         127'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000010000000000000000000000000000000000000000; // D (0x00000000000080000000010000000000) 
14'h2fe5 : LOC =         127'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000010000000000000000000000000000000000000000; // D (0x00000000000100000000010000000000) 
14'h0d87 : LOC =         127'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000010000000000000000000000000000000000000000; // D (0x00000000000200000000010000000000) 
14'h0a34 : LOC =         127'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000010000000000000000000000000000000000000000; // D (0x00000000000400000000010000000000) 
14'h0552 : LOC =         127'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000010000000000000000000000000000000000000000; // D (0x00000000000800000000010000000000) 
14'h1b9e : LOC =         127'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000010000000000000000000000000000000000000000; // D (0x00000000001000000000010000000000) 
14'h2606 : LOC =         127'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000010000000000000000000000000000000000000000; // D (0x00000000002000000000010000000000) 
14'h1e41 : LOC =         127'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000010000000000000000000000000000000000000000; // D (0x00000000004000000000010000000000) 
14'h2db8 : LOC =         127'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000010000000000000000000000000000000000000000; // D (0x00000000008000000000010000000000) 
14'h093d : LOC =         127'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000010000000000000000000000000000000000000000; // D (0x00000000010000000000010000000000) 
14'h0340 : LOC =         127'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000010000000000000000000000000000000000000000; // D (0x00000000020000000000010000000000) 
14'h17ba : LOC =         127'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000; // D (0x00000000040000000000010000000000) 
14'h3e4e : LOC =         127'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000; // D (0x00000000080000000000010000000000) 
14'h2ed1 : LOC =         127'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000; // D (0x00000000100000000000010000000000) 
14'h0fef : LOC =         127'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000; // D (0x00000000200000000000010000000000) 
14'h0ee4 : LOC =         127'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000; // D (0x00000000400000000000010000000000) 
14'h0cf2 : LOC =         127'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000; // D (0x00000000800000000000010000000000) 
14'h08de : LOC =         127'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000; // D (0x00000001000000000000010000000000) 
14'h0086 : LOC =         127'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000; // D (0x00000002000000000000010000000000) 
14'h1036 : LOC =         127'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000; // D (0x00000004000000000000010000000000) 
14'h3156 : LOC =         127'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000; // D (0x00000008000000000000010000000000) 
14'h30e1 : LOC =         127'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000; // D (0x00000010000000000000010000000000) 
14'h338f : LOC =         127'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000; // D (0x00000020000000000000010000000000) 
14'h3553 : LOC =         127'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000; // D (0x00000040000000000000010000000000) 
14'h38eb : LOC =         127'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000; // D (0x00000080000000000000010000000000) 
14'h239b : LOC =         127'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000; // D (0x00000100000000000000010000000000) 
14'h157b : LOC =         127'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000; // D (0x00000200000000000000010000000000) 
14'h3bcc : LOC =         127'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000; // D (0x00000400000000000000010000000000) 
14'h25d5 : LOC =         127'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000; // D (0x00000800000000000000010000000000) 
14'h19e7 : LOC =         127'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000; // D (0x00001000000000000000010000000000) 
14'h22f4 : LOC =         127'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000; // D (0x00002000000000000000010000000000) 
14'h17a5 : LOC =         127'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000; // D (0x00004000000000000000010000000000) 
14'h3e70 : LOC =         127'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000; // D (0x00008000000000000000010000000000) 
14'h2ead : LOC =         127'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000; // D (0x00010000000000000000010000000000) 
14'h0f17 : LOC =         127'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000; // D (0x00020000000000000000010000000000) 
14'h0f14 : LOC =         127'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000; // D (0x00040000000000000000010000000000) 
14'h0f12 : LOC =         127'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000; // D (0x00080000000000000000010000000000) 
14'h0f1e : LOC =         127'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000; // D (0x00100000000000000000010000000000) 
14'h0f06 : LOC =         127'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000; // D (0x00200000000000000000010000000000) 
14'h0f36 : LOC =         127'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000; // D (0x00400000000000000000010000000000) 
14'h0f56 : LOC =         127'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000; // D (0x00800000000000000000010000000000) 
14'h0f96 : LOC =         127'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000; // D (0x01000000000000000000010000000000) 
14'h0e16 : LOC =         127'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000; // D (0x02000000000000000000010000000000) 
14'h0d16 : LOC =         127'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000; // D (0x04000000000000000000010000000000) 
14'h0b16 : LOC =         127'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000; // D (0x08000000000000000000010000000000) 
14'h0716 : LOC =         127'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000; // D (0x10000000000000000000010000000000) 
14'h1f16 : LOC =         127'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000; // D (0x20000000000000000000010000000000) 
14'h2f16 : LOC =         127'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000; // D (0x40000000000000000000010000000000) 
14'h1e2c : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000; // S (0x00000000000000000000020000000000) 
14'h2274 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000000000000000; // D (0x00000000000000000000060000000000) 
14'h25eb : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000000000000000000; // D (0x000000000000000000000a0000000000) 
14'h2ad5 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000; // D (0x00000000000000000000120000000000) 
14'h34a9 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000100000000000000000000000000000000000000000; // D (0x00000000000000000000220000000000) 
14'h0851 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000100000000000000000000000000000000000000000; // D (0x00000000000000000000420000000000) 
14'h32d6 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000100000000000000000000000000000000000000000; // D (0x00000000000000000000820000000000) 
14'h04af : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000100000000000000000000000000000000000000000; // D (0x00000000000000000001020000000000) 
14'h2b2a : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000100000000000000000000000000000000000000000; // D (0x00000000000000000002020000000000) 
14'h3757 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000100000000000000000000000000000000000000000; // D (0x00000000000000000004020000000000) 
14'h0fad : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000100000000000000000000000000000000000000000; // D (0x00000000000000000008020000000000) 
14'h3d2e : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000100000000000000000000000000000000000000000; // D (0x00000000000000000010020000000000) 
14'h1b5f : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000100000000000000000000000000000000000000000; // D (0x00000000000000000020020000000000) 
14'h14ca : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000100000000000000000000000000000000000000000; // D (0x00000000000000000040020000000000) 
14'h0be0 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000100000000000000000000000000000000000000000; // D (0x00000000000000000080020000000000) 
14'h35b4 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000100000000000000000000000000000000000000000; // D (0x00000000000000000100020000000000) 
14'h0a6b : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000100000000000000000000000000000000000000000; // D (0x00000000000000000200020000000000) 
14'h36a2 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000100000000000000000000000000000000000000000; // D (0x00000000000000000400020000000000) 
14'h0c47 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000100000000000000000000000000000000000000000; // D (0x00000000000000000800020000000000) 
14'h3afa : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000100000000000000000000000000000000000000000; // D (0x00000000000000001000020000000000) 
14'h14f7 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000100000000000000000000000000000000000000000; // D (0x00000000000000002000020000000000) 
14'h0b9a : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000100000000000000000000000000000000000000000; // D (0x00000000000000004000020000000000) 
14'h3540 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000100000000000000000000000000000000000000000; // D (0x00000000000000008000020000000000) 
14'h0b83 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000100000000000000000000000000000000000000000; // D (0x00000000000000010000020000000000) 
14'h3572 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000100000000000000000000000000000000000000000; // D (0x00000000000000020000020000000000) 
14'h0be7 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000100000000000000000000000000000000000000000; // D (0x00000000000000040000020000000000) 
14'h35ba : LOC =         127'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000100000000000000000000000000000000000000000; // D (0x00000000000000080000020000000000) 
14'h0a77 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000100000000000000000000000000000000000000000; // D (0x00000000000000100000020000000000) 
14'h369a : LOC =         127'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000100000000000000000000000000000000000000000; // D (0x00000000000000200000020000000000) 
14'h0c37 : LOC =         127'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000100000000000000000000000000000000000000000; // D (0x00000000000000400000020000000000) 
14'h3a1a : LOC =         127'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000100000000000000000000000000000000000000000; // D (0x00000000000000800000020000000000) 
14'h1537 : LOC =         127'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000100000000000000000000000000000000000000000; // D (0x00000000000001000000020000000000) 
14'h081a : LOC =         127'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000100000000000000000000000000000000000000000; // D (0x00000000000002000000020000000000) 
14'h3240 : LOC =         127'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000100000000000000000000000000000000000000000; // D (0x00000000000004000000020000000000) 
14'h0583 : LOC =         127'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000100000000000000000000000000000000000000000; // D (0x00000000000008000000020000000000) 
14'h2972 : LOC =         127'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000100000000000000000000000000000000000000000; // D (0x00000000000010000000020000000000) 
14'h33e7 : LOC =         127'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000100000000000000000000000000000000000000000; // D (0x00000000000020000000020000000000) 
14'h06cd : LOC =         127'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000100000000000000000000000000000000000000000; // D (0x00000000000040000000020000000000) 
14'h2fee : LOC =         127'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000100000000000000000000000000000000000000000; // D (0x00000000000080000000020000000000) 
14'h3edf : LOC =         127'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000100000000000000000000000000000000000000000; // D (0x00000000000100000000020000000000) 
14'h1cbd : LOC =         127'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000100000000000000000000000000000000000000000; // D (0x00000000000200000000020000000000) 
14'h1b0e : LOC =         127'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000100000000000000000000000000000000000000000; // D (0x00000000000400000000020000000000) 
14'h1468 : LOC =         127'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000100000000000000000000000000000000000000000; // D (0x00000000000800000000020000000000) 
14'h0aa4 : LOC =         127'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000100000000000000000000000000000000000000000; // D (0x00000000001000000000020000000000) 
14'h373c : LOC =         127'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000100000000000000000000000000000000000000000; // D (0x00000000002000000000020000000000) 
14'h0f7b : LOC =         127'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000100000000000000000000000000000000000000000; // D (0x00000000004000000000020000000000) 
14'h3c82 : LOC =         127'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000100000000000000000000000000000000000000000; // D (0x00000000008000000000020000000000) 
14'h1807 : LOC =         127'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000100000000000000000000000000000000000000000; // D (0x00000000010000000000020000000000) 
14'h127a : LOC =         127'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000100000000000000000000000000000000000000000; // D (0x00000000020000000000020000000000) 
14'h0680 : LOC =         127'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000; // D (0x00000000040000000000020000000000) 
14'h2f74 : LOC =         127'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000; // D (0x00000000080000000000020000000000) 
14'h3feb : LOC =         127'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000; // D (0x00000000100000000000020000000000) 
14'h1ed5 : LOC =         127'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000; // D (0x00000000200000000000020000000000) 
14'h1fde : LOC =         127'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000; // D (0x00000000400000000000020000000000) 
14'h1dc8 : LOC =         127'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000; // D (0x00000000800000000000020000000000) 
14'h19e4 : LOC =         127'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000; // D (0x00000001000000000000020000000000) 
14'h11bc : LOC =         127'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000; // D (0x00000002000000000000020000000000) 
14'h010c : LOC =         127'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000; // D (0x00000004000000000000020000000000) 
14'h206c : LOC =         127'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000; // D (0x00000008000000000000020000000000) 
14'h21db : LOC =         127'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000; // D (0x00000010000000000000020000000000) 
14'h22b5 : LOC =         127'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000; // D (0x00000020000000000000020000000000) 
14'h2469 : LOC =         127'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000; // D (0x00000040000000000000020000000000) 
14'h29d1 : LOC =         127'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000; // D (0x00000080000000000000020000000000) 
14'h32a1 : LOC =         127'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000; // D (0x00000100000000000000020000000000) 
14'h0441 : LOC =         127'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000; // D (0x00000200000000000000020000000000) 
14'h2af6 : LOC =         127'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000; // D (0x00000400000000000000020000000000) 
14'h34ef : LOC =         127'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000; // D (0x00000800000000000000020000000000) 
14'h08dd : LOC =         127'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000; // D (0x00001000000000000000020000000000) 
14'h33ce : LOC =         127'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000; // D (0x00002000000000000000020000000000) 
14'h069f : LOC =         127'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000; // D (0x00004000000000000000020000000000) 
14'h2f4a : LOC =         127'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000; // D (0x00008000000000000000020000000000) 
14'h3f97 : LOC =         127'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000; // D (0x00010000000000000000020000000000) 
14'h1e2d : LOC =         127'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000; // D (0x00020000000000000000020000000000) 
14'h1e2e : LOC =         127'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000; // D (0x00040000000000000000020000000000) 
14'h1e28 : LOC =         127'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000; // D (0x00080000000000000000020000000000) 
14'h1e24 : LOC =         127'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000; // D (0x00100000000000000000020000000000) 
14'h1e3c : LOC =         127'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000; // D (0x00200000000000000000020000000000) 
14'h1e0c : LOC =         127'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000; // D (0x00400000000000000000020000000000) 
14'h1e6c : LOC =         127'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000; // D (0x00800000000000000000020000000000) 
14'h1eac : LOC =         127'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000; // D (0x01000000000000000000020000000000) 
14'h1f2c : LOC =         127'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000; // D (0x02000000000000000000020000000000) 
14'h1c2c : LOC =         127'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000; // D (0x04000000000000000000020000000000) 
14'h1a2c : LOC =         127'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000; // D (0x08000000000000000000020000000000) 
14'h162c : LOC =         127'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000; // D (0x10000000000000000000020000000000) 
14'h0e2c : LOC =         127'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000; // D (0x20000000000000000000020000000000) 
14'h3e2c : LOC =         127'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000; // D (0x40000000000000000000020000000000) 
14'h3c58 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000; // S (0x00000000000000000000040000000000) 
14'h079f : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000000000000000000000; // D (0x000000000000000000000c0000000000) 
14'h08a1 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000101000000000000000000000000000000000000000000; // D (0x00000000000000000000140000000000) 
14'h16dd : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000; // D (0x00000000000000000000240000000000) 
14'h2a25 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010001000000000000000000000000000000000000000000; // D (0x00000000000000000000440000000000) 
14'h10a2 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100001000000000000000000000000000000000000000000; // D (0x00000000000000000000840000000000) 
14'h26db : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000001000000000000000000000000000000000000000000; // D (0x00000000000000000001040000000000) 
14'h095e : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000001000000000000000000000000000000000000000000; // D (0x00000000000000000002040000000000) 
14'h1523 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000001000000000000000000000000000000000000000000; // D (0x00000000000000000004040000000000) 
14'h2dd9 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000001000000000000000000000000000000000000000000; // D (0x00000000000000000008040000000000) 
14'h1f5a : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000001000000000000000000000000000000000000000000; // D (0x00000000000000000010040000000000) 
14'h392b : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000001000000000000000000000000000000000000000000; // D (0x00000000000000000020040000000000) 
14'h36be : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000001000000000000000000000000000000000000000000; // D (0x00000000000000000040040000000000) 
14'h2994 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000001000000000000000000000000000000000000000000; // D (0x00000000000000000080040000000000) 
14'h17c0 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000001000000000000000000000000000000000000000000; // D (0x00000000000000000100040000000000) 
14'h281f : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000001000000000000000000000000000000000000000000; // D (0x00000000000000000200040000000000) 
14'h14d6 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000001000000000000000000000000000000000000000000; // D (0x00000000000000000400040000000000) 
14'h2e33 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000001000000000000000000000000000000000000000000; // D (0x00000000000000000800040000000000) 
14'h188e : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000001000000000000000000000000000000000000000000; // D (0x00000000000000001000040000000000) 
14'h3683 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000001000000000000000000000000000000000000000000; // D (0x00000000000000002000040000000000) 
14'h29ee : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000001000000000000000000000000000000000000000000; // D (0x00000000000000004000040000000000) 
14'h1734 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000001000000000000000000000000000000000000000000; // D (0x00000000000000008000040000000000) 
14'h29f7 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000001000000000000000000000000000000000000000000; // D (0x00000000000000010000040000000000) 
14'h1706 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000001000000000000000000000000000000000000000000; // D (0x00000000000000020000040000000000) 
14'h2993 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000001000000000000000000000000000000000000000000; // D (0x00000000000000040000040000000000) 
14'h17ce : LOC =         127'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000001000000000000000000000000000000000000000000; // D (0x00000000000000080000040000000000) 
14'h2803 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000001000000000000000000000000000000000000000000; // D (0x00000000000000100000040000000000) 
14'h14ee : LOC =         127'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000001000000000000000000000000000000000000000000; // D (0x00000000000000200000040000000000) 
14'h2e43 : LOC =         127'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000001000000000000000000000000000000000000000000; // D (0x00000000000000400000040000000000) 
14'h186e : LOC =         127'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000001000000000000000000000000000000000000000000; // D (0x00000000000000800000040000000000) 
14'h3743 : LOC =         127'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000001000000000000000000000000000000000000000000; // D (0x00000000000001000000040000000000) 
14'h2a6e : LOC =         127'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000001000000000000000000000000000000000000000000; // D (0x00000000000002000000040000000000) 
14'h1034 : LOC =         127'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000001000000000000000000000000000000000000000000; // D (0x00000000000004000000040000000000) 
14'h27f7 : LOC =         127'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000001000000000000000000000000000000000000000000; // D (0x00000000000008000000040000000000) 
14'h0b06 : LOC =         127'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000000000000000; // D (0x00000000000010000000040000000000) 
14'h1193 : LOC =         127'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000001000000000000000000000000000000000000000000; // D (0x00000000000020000000040000000000) 
14'h24b9 : LOC =         127'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000001000000000000000000000000000000000000000000; // D (0x00000000000040000000040000000000) 
14'h0d9a : LOC =         127'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000001000000000000000000000000000000000000000000; // D (0x00000000000080000000040000000000) 
14'h1cab : LOC =         127'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000000000; // D (0x00000000000100000000040000000000) 
14'h3ec9 : LOC =         127'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000001000000000000000000000000000000000000000000; // D (0x00000000000200000000040000000000) 
14'h397a : LOC =         127'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000001000000000000000000000000000000000000000000; // D (0x00000000000400000000040000000000) 
14'h361c : LOC =         127'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000001000000000000000000000000000000000000000000; // D (0x00000000000800000000040000000000) 
14'h28d0 : LOC =         127'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000001000000000000000000000000000000000000000000; // D (0x00000000001000000000040000000000) 
14'h1548 : LOC =         127'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000001000000000000000000000000000000000000000000; // D (0x00000000002000000000040000000000) 
14'h2d0f : LOC =         127'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000001000000000000000000000000000000000000000000; // D (0x00000000004000000000040000000000) 
14'h1ef6 : LOC =         127'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000001000000000000000000000000000000000000000000; // D (0x00000000008000000000040000000000) 
14'h3a73 : LOC =         127'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000001000000000000000000000000000000000000000000; // D (0x00000000010000000000040000000000) 
14'h300e : LOC =         127'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000001000000000000000000000000000000000000000000; // D (0x00000000020000000000040000000000) 
14'h24f4 : LOC =         127'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000; // D (0x00000000040000000000040000000000) 
14'h0d00 : LOC =         127'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000; // D (0x00000000080000000000040000000000) 
14'h1d9f : LOC =         127'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000; // D (0x00000000100000000000040000000000) 
14'h3ca1 : LOC =         127'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000; // D (0x00000000200000000000040000000000) 
14'h3daa : LOC =         127'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000; // D (0x00000000400000000000040000000000) 
14'h3fbc : LOC =         127'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000; // D (0x00000000800000000000040000000000) 
14'h3b90 : LOC =         127'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000; // D (0x00000001000000000000040000000000) 
14'h33c8 : LOC =         127'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000; // D (0x00000002000000000000040000000000) 
14'h2378 : LOC =         127'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000; // D (0x00000004000000000000040000000000) 
14'h0218 : LOC =         127'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000; // D (0x00000008000000000000040000000000) 
14'h03af : LOC =         127'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000; // D (0x00000010000000000000040000000000) 
14'h00c1 : LOC =         127'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000; // D (0x00000020000000000000040000000000) 
14'h061d : LOC =         127'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000; // D (0x00000040000000000000040000000000) 
14'h0ba5 : LOC =         127'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000; // D (0x00000080000000000000040000000000) 
14'h10d5 : LOC =         127'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000; // D (0x00000100000000000000040000000000) 
14'h2635 : LOC =         127'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000; // D (0x00000200000000000000040000000000) 
14'h0882 : LOC =         127'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000; // D (0x00000400000000000000040000000000) 
14'h169b : LOC =         127'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000; // D (0x00000800000000000000040000000000) 
14'h2aa9 : LOC =         127'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000; // D (0x00001000000000000000040000000000) 
14'h11ba : LOC =         127'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000; // D (0x00002000000000000000040000000000) 
14'h24eb : LOC =         127'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000; // D (0x00004000000000000000040000000000) 
14'h0d3e : LOC =         127'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000; // D (0x00008000000000000000040000000000) 
14'h1de3 : LOC =         127'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000; // D (0x00010000000000000000040000000000) 
14'h3c59 : LOC =         127'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000; // D (0x00020000000000000000040000000000) 
14'h3c5a : LOC =         127'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000; // D (0x00040000000000000000040000000000) 
14'h3c5c : LOC =         127'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000; // D (0x00080000000000000000040000000000) 
14'h3c50 : LOC =         127'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000; // D (0x00100000000000000000040000000000) 
14'h3c48 : LOC =         127'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000; // D (0x00200000000000000000040000000000) 
14'h3c78 : LOC =         127'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000; // D (0x00400000000000000000040000000000) 
14'h3c18 : LOC =         127'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000; // D (0x00800000000000000000040000000000) 
14'h3cd8 : LOC =         127'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000; // D (0x01000000000000000000040000000000) 
14'h3d58 : LOC =         127'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000; // D (0x02000000000000000000040000000000) 
14'h3e58 : LOC =         127'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000; // D (0x04000000000000000000040000000000) 
14'h3858 : LOC =         127'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000; // D (0x08000000000000000000040000000000) 
14'h3458 : LOC =         127'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000; // D (0x10000000000000000000040000000000) 
14'h2c58 : LOC =         127'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000; // D (0x20000000000000000000040000000000) 
14'h1c58 : LOC =         127'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000; // D (0x40000000000000000000040000000000) 
14'h3bc7 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000; // S (0x00000000000000000000080000000000) 
14'h0f3e : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000000000000000000000000; // D (0x00000000000000000000180000000000) 
14'h1142 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001010000000000000000000000000000000000000000000; // D (0x00000000000000000000280000000000) 
14'h2dba : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000; // D (0x00000000000000000000480000000000) 
14'h173d : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100010000000000000000000000000000000000000000000; // D (0x00000000000000000000880000000000) 
14'h2144 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000010000000000000000000000000000000000000000000; // D (0x00000000000000000001080000000000) 
14'h0ec1 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000010000000000000000000000000000000000000000000; // D (0x00000000000000000002080000000000) 
14'h12bc : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000010000000000000000000000000000000000000000000; // D (0x00000000000000000004080000000000) 
14'h2a46 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000010000000000000000000000000000000000000000000; // D (0x00000000000000000008080000000000) 
14'h18c5 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000010000000000000000000000000000000000000000000; // D (0x00000000000000000010080000000000) 
14'h3eb4 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000010000000000000000000000000000000000000000000; // D (0x00000000000000000020080000000000) 
14'h3121 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000010000000000000000000000000000000000000000000; // D (0x00000000000000000040080000000000) 
14'h2e0b : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000010000000000000000000000000000000000000000000; // D (0x00000000000000000080080000000000) 
14'h105f : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000010000000000000000000000000000000000000000000; // D (0x00000000000000000100080000000000) 
14'h2f80 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000010000000000000000000000000000000000000000000; // D (0x00000000000000000200080000000000) 
14'h1349 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000010000000000000000000000000000000000000000000; // D (0x00000000000000000400080000000000) 
14'h29ac : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000010000000000000000000000000000000000000000000; // D (0x00000000000000000800080000000000) 
14'h1f11 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000010000000000000000000000000000000000000000000; // D (0x00000000000000001000080000000000) 
14'h311c : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000010000000000000000000000000000000000000000000; // D (0x00000000000000002000080000000000) 
14'h2e71 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000010000000000000000000000000000000000000000000; // D (0x00000000000000004000080000000000) 
14'h10ab : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000010000000000000000000000000000000000000000000; // D (0x00000000000000008000080000000000) 
14'h2e68 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000010000000000000000000000000000000000000000000; // D (0x00000000000000010000080000000000) 
14'h1099 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000000000000; // D (0x00000000000000020000080000000000) 
14'h2e0c : LOC =         127'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000010000000000000000000000000000000000000000000; // D (0x00000000000000040000080000000000) 
14'h1051 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000010000000000000000000000000000000000000000000; // D (0x00000000000000080000080000000000) 
14'h2f9c : LOC =         127'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000010000000000000000000000000000000000000000000; // D (0x00000000000000100000080000000000) 
14'h1371 : LOC =         127'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000010000000000000000000000000000000000000000000; // D (0x00000000000000200000080000000000) 
14'h29dc : LOC =         127'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000010000000000000000000000000000000000000000000; // D (0x00000000000000400000080000000000) 
14'h1ff1 : LOC =         127'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000010000000000000000000000000000000000000000000; // D (0x00000000000000800000080000000000) 
14'h30dc : LOC =         127'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000010000000000000000000000000000000000000000000; // D (0x00000000000001000000080000000000) 
14'h2df1 : LOC =         127'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000010000000000000000000000000000000000000000000; // D (0x00000000000002000000080000000000) 
14'h17ab : LOC =         127'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000010000000000000000000000000000000000000000000; // D (0x00000000000004000000080000000000) 
14'h2068 : LOC =         127'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000000000000000; // D (0x00000000000008000000080000000000) 
14'h0c99 : LOC =         127'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000010000000000000000000000000000000000000000000; // D (0x00000000000010000000080000000000) 
14'h160c : LOC =         127'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000000000000; // D (0x00000000000020000000080000000000) 
14'h2326 : LOC =         127'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000010000000000000000000000000000000000000000000; // D (0x00000000000040000000080000000000) 
14'h0a05 : LOC =         127'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000010000000000000000000000000000000000000000000; // D (0x00000000000080000000080000000000) 
14'h1b34 : LOC =         127'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000000000000; // D (0x00000000000100000000080000000000) 
14'h3956 : LOC =         127'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000010000000000000000000000000000000000000000000; // D (0x00000000000200000000080000000000) 
14'h3ee5 : LOC =         127'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000010000000000000000000000000000000000000000000; // D (0x00000000000400000000080000000000) 
14'h3183 : LOC =         127'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000010000000000000000000000000000000000000000000; // D (0x00000000000800000000080000000000) 
14'h2f4f : LOC =         127'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000010000000000000000000000000000000000000000000; // D (0x00000000001000000000080000000000) 
14'h12d7 : LOC =         127'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000010000000000000000000000000000000000000000000; // D (0x00000000002000000000080000000000) 
14'h2a90 : LOC =         127'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000010000000000000000000000000000000000000000000; // D (0x00000000004000000000080000000000) 
14'h1969 : LOC =         127'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000010000000000000000000000000000000000000000000; // D (0x00000000008000000000080000000000) 
14'h3dec : LOC =         127'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000010000000000000000000000000000000000000000000; // D (0x00000000010000000000080000000000) 
14'h3791 : LOC =         127'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000010000000000000000000000000000000000000000000; // D (0x00000000020000000000080000000000) 
14'h236b : LOC =         127'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000; // D (0x00000000040000000000080000000000) 
14'h0a9f : LOC =         127'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000; // D (0x00000000080000000000080000000000) 
14'h1a00 : LOC =         127'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000; // D (0x00000000100000000000080000000000) 
14'h3b3e : LOC =         127'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000; // D (0x00000000200000000000080000000000) 
14'h3a35 : LOC =         127'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000; // D (0x00000000400000000000080000000000) 
14'h3823 : LOC =         127'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000; // D (0x00000000800000000000080000000000) 
14'h3c0f : LOC =         127'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000; // D (0x00000001000000000000080000000000) 
14'h3457 : LOC =         127'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000; // D (0x00000002000000000000080000000000) 
14'h24e7 : LOC =         127'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000; // D (0x00000004000000000000080000000000) 
14'h0587 : LOC =         127'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000; // D (0x00000008000000000000080000000000) 
14'h0430 : LOC =         127'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000; // D (0x00000010000000000000080000000000) 
14'h075e : LOC =         127'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000; // D (0x00000020000000000000080000000000) 
14'h0182 : LOC =         127'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000; // D (0x00000040000000000000080000000000) 
14'h0c3a : LOC =         127'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000; // D (0x00000080000000000000080000000000) 
14'h174a : LOC =         127'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000; // D (0x00000100000000000000080000000000) 
14'h21aa : LOC =         127'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000; // D (0x00000200000000000000080000000000) 
14'h0f1d : LOC =         127'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000; // D (0x00000400000000000000080000000000) 
14'h1104 : LOC =         127'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000; // D (0x00000800000000000000080000000000) 
14'h2d36 : LOC =         127'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000; // D (0x00001000000000000000080000000000) 
14'h1625 : LOC =         127'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000; // D (0x00002000000000000000080000000000) 
14'h2374 : LOC =         127'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000; // D (0x00004000000000000000080000000000) 
14'h0aa1 : LOC =         127'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000; // D (0x00008000000000000000080000000000) 
14'h1a7c : LOC =         127'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000; // D (0x00010000000000000000080000000000) 
14'h3bc6 : LOC =         127'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000; // D (0x00020000000000000000080000000000) 
14'h3bc5 : LOC =         127'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000; // D (0x00040000000000000000080000000000) 
14'h3bc3 : LOC =         127'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000; // D (0x00080000000000000000080000000000) 
14'h3bcf : LOC =         127'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000; // D (0x00100000000000000000080000000000) 
14'h3bd7 : LOC =         127'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000; // D (0x00200000000000000000080000000000) 
14'h3be7 : LOC =         127'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000; // D (0x00400000000000000000080000000000) 
14'h3b87 : LOC =         127'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000; // D (0x00800000000000000000080000000000) 
14'h3b47 : LOC =         127'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000; // D (0x01000000000000000000080000000000) 
14'h3ac7 : LOC =         127'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000; // D (0x02000000000000000000080000000000) 
14'h39c7 : LOC =         127'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000; // D (0x04000000000000000000080000000000) 
14'h3fc7 : LOC =         127'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000; // D (0x08000000000000000000080000000000) 
14'h33c7 : LOC =         127'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000; // D (0x10000000000000000000080000000000) 
14'h2bc7 : LOC =         127'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000; // D (0x20000000000000000000080000000000) 
14'h1bc7 : LOC =         127'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000; // D (0x40000000000000000000080000000000) 
14'h34f9 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000; // S (0x00000000000000000000100000000000) 
14'h1e7c : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000000000000000000; // D (0x00000000000000000000300000000000) 
14'h2284 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000000000000000000000; // D (0x00000000000000000000500000000000) 
14'h1803 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000; // D (0x00000000000000000000900000000000) 
14'h2e7a : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000100000000000000000000000000000000000000000000; // D (0x00000000000000000001100000000000) 
14'h01ff : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000100000000000000000000000000000000000000000000; // D (0x00000000000000000002100000000000) 
14'h1d82 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000100000000000000000000000000000000000000000000; // D (0x00000000000000000004100000000000) 
14'h2578 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000100000000000000000000000000000000000000000000; // D (0x00000000000000000008100000000000) 
14'h17fb : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000100000000000000000000000000000000000000000000; // D (0x00000000000000000010100000000000) 
14'h318a : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000100000000000000000000000000000000000000000000; // D (0x00000000000000000020100000000000) 
14'h3e1f : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000100000000000000000000000000000000000000000000; // D (0x00000000000000000040100000000000) 
14'h2135 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000100000000000000000000000000000000000000000000; // D (0x00000000000000000080100000000000) 
14'h1f61 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000100000000000000000000000000000000000000000000; // D (0x00000000000000000100100000000000) 
14'h20be : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000100000000000000000000000000000000000000000000; // D (0x00000000000000000200100000000000) 
14'h1c77 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000100000000000000000000000000000000000000000000; // D (0x00000000000000000400100000000000) 
14'h2692 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000100000000000000000000000000000000000000000000; // D (0x00000000000000000800100000000000) 
14'h102f : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000100000000000000000000000000000000000000000000; // D (0x00000000000000001000100000000000) 
14'h3e22 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000100000000000000000000000000000000000000000000; // D (0x00000000000000002000100000000000) 
14'h214f : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000100000000000000000000000000000000000000000000; // D (0x00000000000000004000100000000000) 
14'h1f95 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000100000000000000000000000000000000000000000000; // D (0x00000000000000008000100000000000) 
14'h2156 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000100000000000000000000000000000000000000000000; // D (0x00000000000000010000100000000000) 
14'h1fa7 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000100000000000000000000000000000000000000000000; // D (0x00000000000000020000100000000000) 
14'h2132 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000100000000000000000000000000000000000000000000; // D (0x00000000000000040000100000000000) 
14'h1f6f : LOC =         127'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000100000000000000000000000000000000000000000000; // D (0x00000000000000080000100000000000) 
14'h20a2 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000100000000000000000000000000000000000000000000; // D (0x00000000000000100000100000000000) 
14'h1c4f : LOC =         127'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000100000000000000000000000000000000000000000000; // D (0x00000000000000200000100000000000) 
14'h26e2 : LOC =         127'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000100000000000000000000000000000000000000000000; // D (0x00000000000000400000100000000000) 
14'h10cf : LOC =         127'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000100000000000000000000000000000000000000000000; // D (0x00000000000000800000100000000000) 
14'h3fe2 : LOC =         127'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000100000000000000000000000000000000000000000000; // D (0x00000000000001000000100000000000) 
14'h22cf : LOC =         127'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000100000000000000000000000000000000000000000000; // D (0x00000000000002000000100000000000) 
14'h1895 : LOC =         127'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000100000000000000000000000000000000000000000000; // D (0x00000000000004000000100000000000) 
14'h2f56 : LOC =         127'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000100000000000000000000000000000000000000000000; // D (0x00000000000008000000100000000000) 
14'h03a7 : LOC =         127'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000100000000000000000000000000000000000000000000; // D (0x00000000000010000000100000000000) 
14'h1932 : LOC =         127'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000100000000000000000000000000000000000000000000; // D (0x00000000000020000000100000000000) 
14'h2c18 : LOC =         127'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000100000000000000000000000000000000000000000000; // D (0x00000000000040000000100000000000) 
14'h053b : LOC =         127'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000100000000000000000000000000000000000000000000; // D (0x00000000000080000000100000000000) 
14'h140a : LOC =         127'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000100000000000000000000000000000000000000000000; // D (0x00000000000100000000100000000000) 
14'h3668 : LOC =         127'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000100000000000000000000000000000000000000000000; // D (0x00000000000200000000100000000000) 
14'h31db : LOC =         127'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000100000000000000000000000000000000000000000000; // D (0x00000000000400000000100000000000) 
14'h3ebd : LOC =         127'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000100000000000000000000000000000000000000000000; // D (0x00000000000800000000100000000000) 
14'h2071 : LOC =         127'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000100000000000000000000000000000000000000000000; // D (0x00000000001000000000100000000000) 
14'h1de9 : LOC =         127'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000100000000000000000000000000000000000000000000; // D (0x00000000002000000000100000000000) 
14'h25ae : LOC =         127'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000100000000000000000000000000000000000000000000; // D (0x00000000004000000000100000000000) 
14'h1657 : LOC =         127'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000100000000000000000000000000000000000000000000; // D (0x00000000008000000000100000000000) 
14'h32d2 : LOC =         127'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000100000000000000000000000000000000000000000000; // D (0x00000000010000000000100000000000) 
14'h38af : LOC =         127'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000100000000000000000000000000000000000000000000; // D (0x00000000020000000000100000000000) 
14'h2c55 : LOC =         127'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000; // D (0x00000000040000000000100000000000) 
14'h05a1 : LOC =         127'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000; // D (0x00000000080000000000100000000000) 
14'h153e : LOC =         127'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000; // D (0x00000000100000000000100000000000) 
14'h3400 : LOC =         127'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000; // D (0x00000000200000000000100000000000) 
14'h350b : LOC =         127'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000; // D (0x00000000400000000000100000000000) 
14'h371d : LOC =         127'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000; // D (0x00000000800000000000100000000000) 
14'h3331 : LOC =         127'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000; // D (0x00000001000000000000100000000000) 
14'h3b69 : LOC =         127'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000; // D (0x00000002000000000000100000000000) 
14'h2bd9 : LOC =         127'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000; // D (0x00000004000000000000100000000000) 
14'h0ab9 : LOC =         127'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000; // D (0x00000008000000000000100000000000) 
14'h0b0e : LOC =         127'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000; // D (0x00000010000000000000100000000000) 
14'h0860 : LOC =         127'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000; // D (0x00000020000000000000100000000000) 
14'h0ebc : LOC =         127'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000; // D (0x00000040000000000000100000000000) 
14'h0304 : LOC =         127'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000; // D (0x00000080000000000000100000000000) 
14'h1874 : LOC =         127'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000; // D (0x00000100000000000000100000000000) 
14'h2e94 : LOC =         127'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000; // D (0x00000200000000000000100000000000) 
14'h0023 : LOC =         127'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000; // D (0x00000400000000000000100000000000) 
14'h1e3a : LOC =         127'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000; // D (0x00000800000000000000100000000000) 
14'h2208 : LOC =         127'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000; // D (0x00001000000000000000100000000000) 
14'h191b : LOC =         127'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000; // D (0x00002000000000000000100000000000) 
14'h2c4a : LOC =         127'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000; // D (0x00004000000000000000100000000000) 
14'h059f : LOC =         127'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000; // D (0x00008000000000000000100000000000) 
14'h1542 : LOC =         127'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000; // D (0x00010000000000000000100000000000) 
14'h34f8 : LOC =         127'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000; // D (0x00020000000000000000100000000000) 
14'h34fb : LOC =         127'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000; // D (0x00040000000000000000100000000000) 
14'h34fd : LOC =         127'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000; // D (0x00080000000000000000100000000000) 
14'h34f1 : LOC =         127'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000; // D (0x00100000000000000000100000000000) 
14'h34e9 : LOC =         127'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000; // D (0x00200000000000000000100000000000) 
14'h34d9 : LOC =         127'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000; // D (0x00400000000000000000100000000000) 
14'h34b9 : LOC =         127'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000; // D (0x00800000000000000000100000000000) 
14'h3479 : LOC =         127'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000; // D (0x01000000000000000000100000000000) 
14'h35f9 : LOC =         127'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000; // D (0x02000000000000000000100000000000) 
14'h36f9 : LOC =         127'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000; // D (0x04000000000000000000100000000000) 
14'h30f9 : LOC =         127'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000; // D (0x08000000000000000000100000000000) 
14'h3cf9 : LOC =         127'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000; // D (0x10000000000000000000100000000000) 
14'h24f9 : LOC =         127'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000; // D (0x20000000000000000000100000000000) 
14'h14f9 : LOC =         127'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000; // D (0x40000000000000000000100000000000) 
14'h2a85 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000; // S (0x00000000000000000000200000000000) 
14'h3cf8 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000000000000000000000000; // D (0x00000000000000000000600000000000) 
14'h067f : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000101000000000000000000000000000000000000000000000; // D (0x00000000000000000000a00000000000) 
14'h3006 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000; // D (0x00000000000000000001200000000000) 
14'h1f83 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000010001000000000000000000000000000000000000000000000; // D (0x00000000000000000002200000000000) 
14'h03fe : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000100001000000000000000000000000000000000000000000000; // D (0x00000000000000000004200000000000) 
14'h3b04 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000001000001000000000000000000000000000000000000000000000; // D (0x00000000000000000008200000000000) 
14'h0987 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000010000001000000000000000000000000000000000000000000000; // D (0x00000000000000000010200000000000) 
14'h2ff6 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000100000001000000000000000000000000000000000000000000000; // D (0x00000000000000000020200000000000) 
14'h2063 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000001000000001000000000000000000000000000000000000000000000; // D (0x00000000000000000040200000000000) 
14'h3f49 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000010000000001000000000000000000000000000000000000000000000; // D (0x00000000000000000080200000000000) 
14'h011d : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000100000000001000000000000000000000000000000000000000000000; // D (0x00000000000000000100200000000000) 
14'h3ec2 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000001000000000001000000000000000000000000000000000000000000000; // D (0x00000000000000000200200000000000) 
14'h020b : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000010000000000001000000000000000000000000000000000000000000000; // D (0x00000000000000000400200000000000) 
14'h38ee : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000100000000000001000000000000000000000000000000000000000000000; // D (0x00000000000000000800200000000000) 
14'h0e53 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000001000000000000001000000000000000000000000000000000000000000000; // D (0x00000000000000001000200000000000) 
14'h205e : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000010000000000000001000000000000000000000000000000000000000000000; // D (0x00000000000000002000200000000000) 
14'h3f33 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000100000000000000001000000000000000000000000000000000000000000000; // D (0x00000000000000004000200000000000) 
14'h01e9 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000001000000000000000001000000000000000000000000000000000000000000000; // D (0x00000000000000008000200000000000) 
14'h3f2a : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000010000000000000000001000000000000000000000000000000000000000000000; // D (0x00000000000000010000200000000000) 
14'h01db : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000100000000000000000001000000000000000000000000000000000000000000000; // D (0x00000000000000020000200000000000) 
14'h3f4e : LOC =         127'b0000000000000000000000000000000000000000000000000000000000001000000000000000000001000000000000000000000000000000000000000000000; // D (0x00000000000000040000200000000000) 
14'h0113 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000010000000000000000000001000000000000000000000000000000000000000000000; // D (0x00000000000000080000200000000000) 
14'h3ede : LOC =         127'b0000000000000000000000000000000000000000000000000000000000100000000000000000000001000000000000000000000000000000000000000000000; // D (0x00000000000000100000200000000000) 
14'h0233 : LOC =         127'b0000000000000000000000000000000000000000000000000000000001000000000000000000000001000000000000000000000000000000000000000000000; // D (0x00000000000000200000200000000000) 
14'h389e : LOC =         127'b0000000000000000000000000000000000000000000000000000000010000000000000000000000001000000000000000000000000000000000000000000000; // D (0x00000000000000400000200000000000) 
14'h0eb3 : LOC =         127'b0000000000000000000000000000000000000000000000000000000100000000000000000000000001000000000000000000000000000000000000000000000; // D (0x00000000000000800000200000000000) 
14'h219e : LOC =         127'b0000000000000000000000000000000000000000000000000000001000000000000000000000000001000000000000000000000000000000000000000000000; // D (0x00000000000001000000200000000000) 
14'h3cb3 : LOC =         127'b0000000000000000000000000000000000000000000000000000010000000000000000000000000001000000000000000000000000000000000000000000000; // D (0x00000000000002000000200000000000) 
14'h06e9 : LOC =         127'b0000000000000000000000000000000000000000000000000000100000000000000000000000000001000000000000000000000000000000000000000000000; // D (0x00000000000004000000200000000000) 
14'h312a : LOC =         127'b0000000000000000000000000000000000000000000000000001000000000000000000000000000001000000000000000000000000000000000000000000000; // D (0x00000000000008000000200000000000) 
14'h1ddb : LOC =         127'b0000000000000000000000000000000000000000000000000010000000000000000000000000000001000000000000000000000000000000000000000000000; // D (0x00000000000010000000200000000000) 
14'h074e : LOC =         127'b0000000000000000000000000000000000000000000000000100000000000000000000000000000001000000000000000000000000000000000000000000000; // D (0x00000000000020000000200000000000) 
14'h3264 : LOC =         127'b0000000000000000000000000000000000000000000000001000000000000000000000000000000001000000000000000000000000000000000000000000000; // D (0x00000000000040000000200000000000) 
14'h1b47 : LOC =         127'b0000000000000000000000000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000000000000000000; // D (0x00000000000080000000200000000000) 
14'h0a76 : LOC =         127'b0000000000000000000000000000000000000000000000100000000000000000000000000000000001000000000000000000000000000000000000000000000; // D (0x00000000000100000000200000000000) 
14'h2814 : LOC =         127'b0000000000000000000000000000000000000000000001000000000000000000000000000000000001000000000000000000000000000000000000000000000; // D (0x00000000000200000000200000000000) 
14'h2fa7 : LOC =         127'b0000000000000000000000000000000000000000000010000000000000000000000000000000000001000000000000000000000000000000000000000000000; // D (0x00000000000400000000200000000000) 
14'h20c1 : LOC =         127'b0000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000000000000; // D (0x00000000000800000000200000000000) 
14'h3e0d : LOC =         127'b0000000000000000000000000000000000000000001000000000000000000000000000000000000001000000000000000000000000000000000000000000000; // D (0x00000000001000000000200000000000) 
14'h0395 : LOC =         127'b0000000000000000000000000000000000000000010000000000000000000000000000000000000001000000000000000000000000000000000000000000000; // D (0x00000000002000000000200000000000) 
14'h3bd2 : LOC =         127'b0000000000000000000000000000000000000000100000000000000000000000000000000000000001000000000000000000000000000000000000000000000; // D (0x00000000004000000000200000000000) 
14'h082b : LOC =         127'b0000000000000000000000000000000000000001000000000000000000000000000000000000000001000000000000000000000000000000000000000000000; // D (0x00000000008000000000200000000000) 
14'h2cae : LOC =         127'b0000000000000000000000000000000000000010000000000000000000000000000000000000000001000000000000000000000000000000000000000000000; // D (0x00000000010000000000200000000000) 
14'h26d3 : LOC =         127'b0000000000000000000000000000000000000100000000000000000000000000000000000000000001000000000000000000000000000000000000000000000; // D (0x00000000020000000000200000000000) 
14'h3229 : LOC =         127'b0000000000000000000000000000000000001000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000; // D (0x00000000040000000000200000000000) 
14'h1bdd : LOC =         127'b0000000000000000000000000000000000010000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000; // D (0x00000000080000000000200000000000) 
14'h0b42 : LOC =         127'b0000000000000000000000000000000000100000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000; // D (0x00000000100000000000200000000000) 
14'h2a7c : LOC =         127'b0000000000000000000000000000000001000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000; // D (0x00000000200000000000200000000000) 
14'h2b77 : LOC =         127'b0000000000000000000000000000000010000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000; // D (0x00000000400000000000200000000000) 
14'h2961 : LOC =         127'b0000000000000000000000000000000100000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000; // D (0x00000000800000000000200000000000) 
14'h2d4d : LOC =         127'b0000000000000000000000000000001000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000; // D (0x00000001000000000000200000000000) 
14'h2515 : LOC =         127'b0000000000000000000000000000010000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000; // D (0x00000002000000000000200000000000) 
14'h35a5 : LOC =         127'b0000000000000000000000000000100000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000; // D (0x00000004000000000000200000000000) 
14'h14c5 : LOC =         127'b0000000000000000000000000001000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000; // D (0x00000008000000000000200000000000) 
14'h1572 : LOC =         127'b0000000000000000000000000010000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000; // D (0x00000010000000000000200000000000) 
14'h161c : LOC =         127'b0000000000000000000000000100000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000; // D (0x00000020000000000000200000000000) 
14'h10c0 : LOC =         127'b0000000000000000000000001000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000; // D (0x00000040000000000000200000000000) 
14'h1d78 : LOC =         127'b0000000000000000000000010000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000; // D (0x00000080000000000000200000000000) 
14'h0608 : LOC =         127'b0000000000000000000000100000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000; // D (0x00000100000000000000200000000000) 
14'h30e8 : LOC =         127'b0000000000000000000001000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000; // D (0x00000200000000000000200000000000) 
14'h1e5f : LOC =         127'b0000000000000000000010000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000; // D (0x00000400000000000000200000000000) 
14'h0046 : LOC =         127'b0000000000000000000100000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000; // D (0x00000800000000000000200000000000) 
14'h3c74 : LOC =         127'b0000000000000000001000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000; // D (0x00001000000000000000200000000000) 
14'h0767 : LOC =         127'b0000000000000000010000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000; // D (0x00002000000000000000200000000000) 
14'h3236 : LOC =         127'b0000000000000000100000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000; // D (0x00004000000000000000200000000000) 
14'h1be3 : LOC =         127'b0000000000000001000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000; // D (0x00008000000000000000200000000000) 
14'h0b3e : LOC =         127'b0000000000000010000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000; // D (0x00010000000000000000200000000000) 
14'h2a84 : LOC =         127'b0000000000000100000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000; // D (0x00020000000000000000200000000000) 
14'h2a87 : LOC =         127'b0000000000001000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000; // D (0x00040000000000000000200000000000) 
14'h2a81 : LOC =         127'b0000000000010000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000; // D (0x00080000000000000000200000000000) 
14'h2a8d : LOC =         127'b0000000000100000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000; // D (0x00100000000000000000200000000000) 
14'h2a95 : LOC =         127'b0000000001000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000; // D (0x00200000000000000000200000000000) 
14'h2aa5 : LOC =         127'b0000000010000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000; // D (0x00400000000000000000200000000000) 
14'h2ac5 : LOC =         127'b0000000100000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000; // D (0x00800000000000000000200000000000) 
14'h2a05 : LOC =         127'b0000001000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000; // D (0x01000000000000000000200000000000) 
14'h2b85 : LOC =         127'b0000010000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000; // D (0x02000000000000000000200000000000) 
14'h2885 : LOC =         127'b0000100000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000; // D (0x04000000000000000000200000000000) 
14'h2e85 : LOC =         127'b0001000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000; // D (0x08000000000000000000200000000000) 
14'h2285 : LOC =         127'b0010000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000; // D (0x10000000000000000000200000000000) 
14'h3a85 : LOC =         127'b0100000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000; // D (0x20000000000000000000200000000000) 
14'h0a85 : LOC =         127'b1000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000; // D (0x40000000000000000000200000000000) 
14'h167d : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000; // S (0x00000000000000000000400000000000) 
14'h3a87 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000000000000000000000000000; // D (0x00000000000000000000c00000000000) 
14'h0cfe : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000001010000000000000000000000000000000000000000000000; // D (0x00000000000000000001400000000000) 
14'h237b : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000; // D (0x00000000000000000002400000000000) 
14'h3f06 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000100010000000000000000000000000000000000000000000000; // D (0x00000000000000000004400000000000) 
14'h07fc : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000001000010000000000000000000000000000000000000000000000; // D (0x00000000000000000008400000000000) 
14'h357f : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000010000010000000000000000000000000000000000000000000000; // D (0x00000000000000000010400000000000) 
14'h130e : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000100000010000000000000000000000000000000000000000000000; // D (0x00000000000000000020400000000000) 
14'h1c9b : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000001000000010000000000000000000000000000000000000000000000; // D (0x00000000000000000040400000000000) 
14'h03b1 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000010000000010000000000000000000000000000000000000000000000; // D (0x00000000000000000080400000000000) 
14'h3de5 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000100000000010000000000000000000000000000000000000000000000; // D (0x00000000000000000100400000000000) 
14'h023a : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000001000000000010000000000000000000000000000000000000000000000; // D (0x00000000000000000200400000000000) 
14'h3ef3 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000010000000000010000000000000000000000000000000000000000000000; // D (0x00000000000000000400400000000000) 
14'h0416 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000100000000000010000000000000000000000000000000000000000000000; // D (0x00000000000000000800400000000000) 
14'h32ab : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000001000000000000010000000000000000000000000000000000000000000000; // D (0x00000000000000001000400000000000) 
14'h1ca6 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000010000000000000010000000000000000000000000000000000000000000000; // D (0x00000000000000002000400000000000) 
14'h03cb : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000100000000000000010000000000000000000000000000000000000000000000; // D (0x00000000000000004000400000000000) 
14'h3d11 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000001000000000000000010000000000000000000000000000000000000000000000; // D (0x00000000000000008000400000000000) 
14'h03d2 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000010000000000000000010000000000000000000000000000000000000000000000; // D (0x00000000000000010000400000000000) 
14'h3d23 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000100000000000000000010000000000000000000000000000000000000000000000; // D (0x00000000000000020000400000000000) 
14'h03b6 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000001000000000000000000010000000000000000000000000000000000000000000000; // D (0x00000000000000040000400000000000) 
14'h3deb : LOC =         127'b0000000000000000000000000000000000000000000000000000000000010000000000000000000010000000000000000000000000000000000000000000000; // D (0x00000000000000080000400000000000) 
14'h0226 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000000000000000; // D (0x00000000000000100000400000000000) 
14'h3ecb : LOC =         127'b0000000000000000000000000000000000000000000000000000000001000000000000000000000010000000000000000000000000000000000000000000000; // D (0x00000000000000200000400000000000) 
14'h0466 : LOC =         127'b0000000000000000000000000000000000000000000000000000000010000000000000000000000010000000000000000000000000000000000000000000000; // D (0x00000000000000400000400000000000) 
14'h324b : LOC =         127'b0000000000000000000000000000000000000000000000000000000100000000000000000000000010000000000000000000000000000000000000000000000; // D (0x00000000000000800000400000000000) 
14'h1d66 : LOC =         127'b0000000000000000000000000000000000000000000000000000001000000000000000000000000010000000000000000000000000000000000000000000000; // D (0x00000000000001000000400000000000) 
14'h004b : LOC =         127'b0000000000000000000000000000000000000000000000000000010000000000000000000000000010000000000000000000000000000000000000000000000; // D (0x00000000000002000000400000000000) 
14'h3a11 : LOC =         127'b0000000000000000000000000000000000000000000000000000100000000000000000000000000010000000000000000000000000000000000000000000000; // D (0x00000000000004000000400000000000) 
14'h0dd2 : LOC =         127'b0000000000000000000000000000000000000000000000000001000000000000000000000000000010000000000000000000000000000000000000000000000; // D (0x00000000000008000000400000000000) 
14'h2123 : LOC =         127'b0000000000000000000000000000000000000000000000000010000000000000000000000000000010000000000000000000000000000000000000000000000; // D (0x00000000000010000000400000000000) 
14'h3bb6 : LOC =         127'b0000000000000000000000000000000000000000000000000100000000000000000000000000000010000000000000000000000000000000000000000000000; // D (0x00000000000020000000400000000000) 
14'h0e9c : LOC =         127'b0000000000000000000000000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000000000000000000; // D (0x00000000000040000000400000000000) 
14'h27bf : LOC =         127'b0000000000000000000000000000000000000000000000010000000000000000000000000000000010000000000000000000000000000000000000000000000; // D (0x00000000000080000000400000000000) 
14'h368e : LOC =         127'b0000000000000000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000000000000000; // D (0x00000000000100000000400000000000) 
14'h14ec : LOC =         127'b0000000000000000000000000000000000000000000001000000000000000000000000000000000010000000000000000000000000000000000000000000000; // D (0x00000000000200000000400000000000) 
14'h135f : LOC =         127'b0000000000000000000000000000000000000000000010000000000000000000000000000000000010000000000000000000000000000000000000000000000; // D (0x00000000000400000000400000000000) 
14'h1c39 : LOC =         127'b0000000000000000000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000000000000000; // D (0x00000000000800000000400000000000) 
14'h02f5 : LOC =         127'b0000000000000000000000000000000000000000001000000000000000000000000000000000000010000000000000000000000000000000000000000000000; // D (0x00000000001000000000400000000000) 
14'h3f6d : LOC =         127'b0000000000000000000000000000000000000000010000000000000000000000000000000000000010000000000000000000000000000000000000000000000; // D (0x00000000002000000000400000000000) 
14'h072a : LOC =         127'b0000000000000000000000000000000000000000100000000000000000000000000000000000000010000000000000000000000000000000000000000000000; // D (0x00000000004000000000400000000000) 
14'h34d3 : LOC =         127'b0000000000000000000000000000000000000001000000000000000000000000000000000000000010000000000000000000000000000000000000000000000; // D (0x00000000008000000000400000000000) 
14'h1056 : LOC =         127'b0000000000000000000000000000000000000010000000000000000000000000000000000000000010000000000000000000000000000000000000000000000; // D (0x00000000010000000000400000000000) 
14'h1a2b : LOC =         127'b0000000000000000000000000000000000000100000000000000000000000000000000000000000010000000000000000000000000000000000000000000000; // D (0x00000000020000000000400000000000) 
14'h0ed1 : LOC =         127'b0000000000000000000000000000000000001000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000; // D (0x00000000040000000000400000000000) 
14'h2725 : LOC =         127'b0000000000000000000000000000000000010000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000; // D (0x00000000080000000000400000000000) 
14'h37ba : LOC =         127'b0000000000000000000000000000000000100000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000; // D (0x00000000100000000000400000000000) 
14'h1684 : LOC =         127'b0000000000000000000000000000000001000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000; // D (0x00000000200000000000400000000000) 
14'h178f : LOC =         127'b0000000000000000000000000000000010000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000; // D (0x00000000400000000000400000000000) 
14'h1599 : LOC =         127'b0000000000000000000000000000000100000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000; // D (0x00000000800000000000400000000000) 
14'h11b5 : LOC =         127'b0000000000000000000000000000001000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000; // D (0x00000001000000000000400000000000) 
14'h19ed : LOC =         127'b0000000000000000000000000000010000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000; // D (0x00000002000000000000400000000000) 
14'h095d : LOC =         127'b0000000000000000000000000000100000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000; // D (0x00000004000000000000400000000000) 
14'h283d : LOC =         127'b0000000000000000000000000001000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000; // D (0x00000008000000000000400000000000) 
14'h298a : LOC =         127'b0000000000000000000000000010000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000; // D (0x00000010000000000000400000000000) 
14'h2ae4 : LOC =         127'b0000000000000000000000000100000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000; // D (0x00000020000000000000400000000000) 
14'h2c38 : LOC =         127'b0000000000000000000000001000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000; // D (0x00000040000000000000400000000000) 
14'h2180 : LOC =         127'b0000000000000000000000010000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000; // D (0x00000080000000000000400000000000) 
14'h3af0 : LOC =         127'b0000000000000000000000100000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000; // D (0x00000100000000000000400000000000) 
14'h0c10 : LOC =         127'b0000000000000000000001000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000; // D (0x00000200000000000000400000000000) 
14'h22a7 : LOC =         127'b0000000000000000000010000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000; // D (0x00000400000000000000400000000000) 
14'h3cbe : LOC =         127'b0000000000000000000100000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000; // D (0x00000800000000000000400000000000) 
14'h008c : LOC =         127'b0000000000000000001000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000; // D (0x00001000000000000000400000000000) 
14'h3b9f : LOC =         127'b0000000000000000010000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000; // D (0x00002000000000000000400000000000) 
14'h0ece : LOC =         127'b0000000000000000100000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000; // D (0x00004000000000000000400000000000) 
14'h271b : LOC =         127'b0000000000000001000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000; // D (0x00008000000000000000400000000000) 
14'h37c6 : LOC =         127'b0000000000000010000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000; // D (0x00010000000000000000400000000000) 
14'h167c : LOC =         127'b0000000000000100000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000; // D (0x00020000000000000000400000000000) 
14'h167f : LOC =         127'b0000000000001000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000; // D (0x00040000000000000000400000000000) 
14'h1679 : LOC =         127'b0000000000010000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000; // D (0x00080000000000000000400000000000) 
14'h1675 : LOC =         127'b0000000000100000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000; // D (0x00100000000000000000400000000000) 
14'h166d : LOC =         127'b0000000001000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000; // D (0x00200000000000000000400000000000) 
14'h165d : LOC =         127'b0000000010000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000; // D (0x00400000000000000000400000000000) 
14'h163d : LOC =         127'b0000000100000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000; // D (0x00800000000000000000400000000000) 
14'h16fd : LOC =         127'b0000001000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000; // D (0x01000000000000000000400000000000) 
14'h177d : LOC =         127'b0000010000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000; // D (0x02000000000000000000400000000000) 
14'h147d : LOC =         127'b0000100000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000; // D (0x04000000000000000000400000000000) 
14'h127d : LOC =         127'b0001000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000; // D (0x08000000000000000000400000000000) 
14'h1e7d : LOC =         127'b0010000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000; // D (0x10000000000000000000400000000000) 
14'h067d : LOC =         127'b0100000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000; // D (0x20000000000000000000400000000000) 
14'h367d : LOC =         127'b1000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000; // D (0x40000000000000000000400000000000) 
14'h2cfa : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000; // S (0x00000000000000000000800000000000) 
14'h3679 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000000000000000000000; // D (0x00000000000000000001800000000000) 
14'h19fc : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000000000000000000000000; // D (0x00000000000000000002800000000000) 
14'h0581 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000; // D (0x00000000000000000004800000000000) 
14'h3d7b : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000001000100000000000000000000000000000000000000000000000; // D (0x00000000000000000008800000000000) 
14'h0ff8 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000010000100000000000000000000000000000000000000000000000; // D (0x00000000000000000010800000000000) 
14'h2989 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000100000100000000000000000000000000000000000000000000000; // D (0x00000000000000000020800000000000) 
14'h261c : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000001000000100000000000000000000000000000000000000000000000; // D (0x00000000000000000040800000000000) 
14'h3936 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000010000000100000000000000000000000000000000000000000000000; // D (0x00000000000000000080800000000000) 
14'h0762 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000100000000100000000000000000000000000000000000000000000000; // D (0x00000000000000000100800000000000) 
14'h38bd : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000001000000000100000000000000000000000000000000000000000000000; // D (0x00000000000000000200800000000000) 
14'h0474 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000010000000000100000000000000000000000000000000000000000000000; // D (0x00000000000000000400800000000000) 
14'h3e91 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000100000000000100000000000000000000000000000000000000000000000; // D (0x00000000000000000800800000000000) 
14'h082c : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000001000000000000100000000000000000000000000000000000000000000000; // D (0x00000000000000001000800000000000) 
14'h2621 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000010000000000000100000000000000000000000000000000000000000000000; // D (0x00000000000000002000800000000000) 
14'h394c : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000100000000000000100000000000000000000000000000000000000000000000; // D (0x00000000000000004000800000000000) 
14'h0796 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000001000000000000000100000000000000000000000000000000000000000000000; // D (0x00000000000000008000800000000000) 
14'h3955 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000010000000000000000100000000000000000000000000000000000000000000000; // D (0x00000000000000010000800000000000) 
14'h07a4 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000100000000000000000100000000000000000000000000000000000000000000000; // D (0x00000000000000020000800000000000) 
14'h3931 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000001000000000000000000100000000000000000000000000000000000000000000000; // D (0x00000000000000040000800000000000) 
14'h076c : LOC =         127'b0000000000000000000000000000000000000000000000000000000000010000000000000000000100000000000000000000000000000000000000000000000; // D (0x00000000000000080000800000000000) 
14'h38a1 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000100000000000000000000100000000000000000000000000000000000000000000000; // D (0x00000000000000100000800000000000) 
14'h044c : LOC =         127'b0000000000000000000000000000000000000000000000000000000001000000000000000000000100000000000000000000000000000000000000000000000; // D (0x00000000000000200000800000000000) 
14'h3ee1 : LOC =         127'b0000000000000000000000000000000000000000000000000000000010000000000000000000000100000000000000000000000000000000000000000000000; // D (0x00000000000000400000800000000000) 
14'h08cc : LOC =         127'b0000000000000000000000000000000000000000000000000000000100000000000000000000000100000000000000000000000000000000000000000000000; // D (0x00000000000000800000800000000000) 
14'h27e1 : LOC =         127'b0000000000000000000000000000000000000000000000000000001000000000000000000000000100000000000000000000000000000000000000000000000; // D (0x00000000000001000000800000000000) 
14'h3acc : LOC =         127'b0000000000000000000000000000000000000000000000000000010000000000000000000000000100000000000000000000000000000000000000000000000; // D (0x00000000000002000000800000000000) 
14'h0096 : LOC =         127'b0000000000000000000000000000000000000000000000000000100000000000000000000000000100000000000000000000000000000000000000000000000; // D (0x00000000000004000000800000000000) 
14'h3755 : LOC =         127'b0000000000000000000000000000000000000000000000000001000000000000000000000000000100000000000000000000000000000000000000000000000; // D (0x00000000000008000000800000000000) 
14'h1ba4 : LOC =         127'b0000000000000000000000000000000000000000000000000010000000000000000000000000000100000000000000000000000000000000000000000000000; // D (0x00000000000010000000800000000000) 
14'h0131 : LOC =         127'b0000000000000000000000000000000000000000000000000100000000000000000000000000000100000000000000000000000000000000000000000000000; // D (0x00000000000020000000800000000000) 
14'h341b : LOC =         127'b0000000000000000000000000000000000000000000000001000000000000000000000000000000100000000000000000000000000000000000000000000000; // D (0x00000000000040000000800000000000) 
14'h1d38 : LOC =         127'b0000000000000000000000000000000000000000000000010000000000000000000000000000000100000000000000000000000000000000000000000000000; // D (0x00000000000080000000800000000000) 
14'h0c09 : LOC =         127'b0000000000000000000000000000000000000000000000100000000000000000000000000000000100000000000000000000000000000000000000000000000; // D (0x00000000000100000000800000000000) 
14'h2e6b : LOC =         127'b0000000000000000000000000000000000000000000001000000000000000000000000000000000100000000000000000000000000000000000000000000000; // D (0x00000000000200000000800000000000) 
14'h29d8 : LOC =         127'b0000000000000000000000000000000000000000000010000000000000000000000000000000000100000000000000000000000000000000000000000000000; // D (0x00000000000400000000800000000000) 
14'h26be : LOC =         127'b0000000000000000000000000000000000000000000100000000000000000000000000000000000100000000000000000000000000000000000000000000000; // D (0x00000000000800000000800000000000) 
14'h3872 : LOC =         127'b0000000000000000000000000000000000000000001000000000000000000000000000000000000100000000000000000000000000000000000000000000000; // D (0x00000000001000000000800000000000) 
14'h05ea : LOC =         127'b0000000000000000000000000000000000000000010000000000000000000000000000000000000100000000000000000000000000000000000000000000000; // D (0x00000000002000000000800000000000) 
14'h3dad : LOC =         127'b0000000000000000000000000000000000000000100000000000000000000000000000000000000100000000000000000000000000000000000000000000000; // D (0x00000000004000000000800000000000) 
14'h0e54 : LOC =         127'b0000000000000000000000000000000000000001000000000000000000000000000000000000000100000000000000000000000000000000000000000000000; // D (0x00000000008000000000800000000000) 
14'h2ad1 : LOC =         127'b0000000000000000000000000000000000000010000000000000000000000000000000000000000100000000000000000000000000000000000000000000000; // D (0x00000000010000000000800000000000) 
14'h20ac : LOC =         127'b0000000000000000000000000000000000000100000000000000000000000000000000000000000100000000000000000000000000000000000000000000000; // D (0x00000000020000000000800000000000) 
14'h3456 : LOC =         127'b0000000000000000000000000000000000001000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000; // D (0x00000000040000000000800000000000) 
14'h1da2 : LOC =         127'b0000000000000000000000000000000000010000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000; // D (0x00000000080000000000800000000000) 
14'h0d3d : LOC =         127'b0000000000000000000000000000000000100000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000; // D (0x00000000100000000000800000000000) 
14'h2c03 : LOC =         127'b0000000000000000000000000000000001000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000; // D (0x00000000200000000000800000000000) 
14'h2d08 : LOC =         127'b0000000000000000000000000000000010000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000; // D (0x00000000400000000000800000000000) 
14'h2f1e : LOC =         127'b0000000000000000000000000000000100000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000; // D (0x00000000800000000000800000000000) 
14'h2b32 : LOC =         127'b0000000000000000000000000000001000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000; // D (0x00000001000000000000800000000000) 
14'h236a : LOC =         127'b0000000000000000000000000000010000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000; // D (0x00000002000000000000800000000000) 
14'h33da : LOC =         127'b0000000000000000000000000000100000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000; // D (0x00000004000000000000800000000000) 
14'h12ba : LOC =         127'b0000000000000000000000000001000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000; // D (0x00000008000000000000800000000000) 
14'h130d : LOC =         127'b0000000000000000000000000010000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000; // D (0x00000010000000000000800000000000) 
14'h1063 : LOC =         127'b0000000000000000000000000100000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000; // D (0x00000020000000000000800000000000) 
14'h16bf : LOC =         127'b0000000000000000000000001000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000; // D (0x00000040000000000000800000000000) 
14'h1b07 : LOC =         127'b0000000000000000000000010000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000; // D (0x00000080000000000000800000000000) 
14'h0077 : LOC =         127'b0000000000000000000000100000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000; // D (0x00000100000000000000800000000000) 
14'h3697 : LOC =         127'b0000000000000000000001000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000; // D (0x00000200000000000000800000000000) 
14'h1820 : LOC =         127'b0000000000000000000010000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000; // D (0x00000400000000000000800000000000) 
14'h0639 : LOC =         127'b0000000000000000000100000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000; // D (0x00000800000000000000800000000000) 
14'h3a0b : LOC =         127'b0000000000000000001000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000; // D (0x00001000000000000000800000000000) 
14'h0118 : LOC =         127'b0000000000000000010000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000; // D (0x00002000000000000000800000000000) 
14'h3449 : LOC =         127'b0000000000000000100000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000; // D (0x00004000000000000000800000000000) 
14'h1d9c : LOC =         127'b0000000000000001000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000; // D (0x00008000000000000000800000000000) 
14'h0d41 : LOC =         127'b0000000000000010000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000; // D (0x00010000000000000000800000000000) 
14'h2cfb : LOC =         127'b0000000000000100000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000; // D (0x00020000000000000000800000000000) 
14'h2cf8 : LOC =         127'b0000000000001000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000; // D (0x00040000000000000000800000000000) 
14'h2cfe : LOC =         127'b0000000000010000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000; // D (0x00080000000000000000800000000000) 
14'h2cf2 : LOC =         127'b0000000000100000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000; // D (0x00100000000000000000800000000000) 
14'h2cea : LOC =         127'b0000000001000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000; // D (0x00200000000000000000800000000000) 
14'h2cda : LOC =         127'b0000000010000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000; // D (0x00400000000000000000800000000000) 
14'h2cba : LOC =         127'b0000000100000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000; // D (0x00800000000000000000800000000000) 
14'h2c7a : LOC =         127'b0000001000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000; // D (0x01000000000000000000800000000000) 
14'h2dfa : LOC =         127'b0000010000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000; // D (0x02000000000000000000800000000000) 
14'h2efa : LOC =         127'b0000100000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000; // D (0x04000000000000000000800000000000) 
14'h28fa : LOC =         127'b0001000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000; // D (0x08000000000000000000800000000000) 
14'h24fa : LOC =         127'b0010000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000; // D (0x10000000000000000000800000000000) 
14'h3cfa : LOC =         127'b0100000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000; // D (0x20000000000000000000800000000000) 
14'h0cfa : LOC =         127'b1000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000; // D (0x40000000000000000000800000000000) 
14'h1a83 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000; // S (0x00000000000000000001000000000000) 
14'h2f85 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000000000000000000000000000; // D (0x00000000000000000003000000000000) 
14'h33f8 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000101000000000000000000000000000000000000000000000000; // D (0x00000000000000000005000000000000) 
14'h0b02 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000; // D (0x00000000000000000009000000000000) 
14'h3981 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000010001000000000000000000000000000000000000000000000000; // D (0x00000000000000000011000000000000) 
14'h1ff0 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000100001000000000000000000000000000000000000000000000000; // D (0x00000000000000000021000000000000) 
14'h1065 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000001000001000000000000000000000000000000000000000000000000; // D (0x00000000000000000041000000000000) 
14'h0f4f : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000010000001000000000000000000000000000000000000000000000000; // D (0x00000000000000000081000000000000) 
14'h311b : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000100000001000000000000000000000000000000000000000000000000; // D (0x00000000000000000101000000000000) 
14'h0ec4 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000001000000001000000000000000000000000000000000000000000000000; // D (0x00000000000000000201000000000000) 
14'h320d : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000010000000001000000000000000000000000000000000000000000000000; // D (0x00000000000000000401000000000000) 
14'h08e8 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000100000000001000000000000000000000000000000000000000000000000; // D (0x00000000000000000801000000000000) 
14'h3e55 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000001000000000001000000000000000000000000000000000000000000000000; // D (0x00000000000000001001000000000000) 
14'h1058 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000010000000000001000000000000000000000000000000000000000000000000; // D (0x00000000000000002001000000000000) 
14'h0f35 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000100000000000001000000000000000000000000000000000000000000000000; // D (0x00000000000000004001000000000000) 
14'h31ef : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000001000000000000001000000000000000000000000000000000000000000000000; // D (0x00000000000000008001000000000000) 
14'h0f2c : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000010000000000000001000000000000000000000000000000000000000000000000; // D (0x00000000000000010001000000000000) 
14'h31dd : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000100000000000000001000000000000000000000000000000000000000000000000; // D (0x00000000000000020001000000000000) 
14'h0f48 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000001000000000000000001000000000000000000000000000000000000000000000000; // D (0x00000000000000040001000000000000) 
14'h3115 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000010000000000000000001000000000000000000000000000000000000000000000000; // D (0x00000000000000080001000000000000) 
14'h0ed8 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000100000000000000000001000000000000000000000000000000000000000000000000; // D (0x00000000000000100001000000000000) 
14'h3235 : LOC =         127'b0000000000000000000000000000000000000000000000000000000001000000000000000000001000000000000000000000000000000000000000000000000; // D (0x00000000000000200001000000000000) 
14'h0898 : LOC =         127'b0000000000000000000000000000000000000000000000000000000010000000000000000000001000000000000000000000000000000000000000000000000; // D (0x00000000000000400001000000000000) 
14'h3eb5 : LOC =         127'b0000000000000000000000000000000000000000000000000000000100000000000000000000001000000000000000000000000000000000000000000000000; // D (0x00000000000000800001000000000000) 
14'h1198 : LOC =         127'b0000000000000000000000000000000000000000000000000000001000000000000000000000001000000000000000000000000000000000000000000000000; // D (0x00000000000001000001000000000000) 
14'h0cb5 : LOC =         127'b0000000000000000000000000000000000000000000000000000010000000000000000000000001000000000000000000000000000000000000000000000000; // D (0x00000000000002000001000000000000) 
14'h36ef : LOC =         127'b0000000000000000000000000000000000000000000000000000100000000000000000000000001000000000000000000000000000000000000000000000000; // D (0x00000000000004000001000000000000) 
14'h012c : LOC =         127'b0000000000000000000000000000000000000000000000000001000000000000000000000000001000000000000000000000000000000000000000000000000; // D (0x00000000000008000001000000000000) 
14'h2ddd : LOC =         127'b0000000000000000000000000000000000000000000000000010000000000000000000000000001000000000000000000000000000000000000000000000000; // D (0x00000000000010000001000000000000) 
14'h3748 : LOC =         127'b0000000000000000000000000000000000000000000000000100000000000000000000000000001000000000000000000000000000000000000000000000000; // D (0x00000000000020000001000000000000) 
14'h0262 : LOC =         127'b0000000000000000000000000000000000000000000000001000000000000000000000000000001000000000000000000000000000000000000000000000000; // D (0x00000000000040000001000000000000) 
14'h2b41 : LOC =         127'b0000000000000000000000000000000000000000000000010000000000000000000000000000001000000000000000000000000000000000000000000000000; // D (0x00000000000080000001000000000000) 
14'h3a70 : LOC =         127'b0000000000000000000000000000000000000000000000100000000000000000000000000000001000000000000000000000000000000000000000000000000; // D (0x00000000000100000001000000000000) 
14'h1812 : LOC =         127'b0000000000000000000000000000000000000000000001000000000000000000000000000000001000000000000000000000000000000000000000000000000; // D (0x00000000000200000001000000000000) 
14'h1fa1 : LOC =         127'b0000000000000000000000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000000000000000000000; // D (0x00000000000400000001000000000000) 
14'h10c7 : LOC =         127'b0000000000000000000000000000000000000000000100000000000000000000000000000000001000000000000000000000000000000000000000000000000; // D (0x00000000000800000001000000000000) 
14'h0e0b : LOC =         127'b0000000000000000000000000000000000000000001000000000000000000000000000000000001000000000000000000000000000000000000000000000000; // D (0x00000000001000000001000000000000) 
14'h3393 : LOC =         127'b0000000000000000000000000000000000000000010000000000000000000000000000000000001000000000000000000000000000000000000000000000000; // D (0x00000000002000000001000000000000) 
14'h0bd4 : LOC =         127'b0000000000000000000000000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000000000000000; // D (0x00000000004000000001000000000000) 
14'h382d : LOC =         127'b0000000000000000000000000000000000000001000000000000000000000000000000000000001000000000000000000000000000000000000000000000000; // D (0x00000000008000000001000000000000) 
14'h1ca8 : LOC =         127'b0000000000000000000000000000000000000010000000000000000000000000000000000000001000000000000000000000000000000000000000000000000; // D (0x00000000010000000001000000000000) 
14'h16d5 : LOC =         127'b0000000000000000000000000000000000000100000000000000000000000000000000000000001000000000000000000000000000000000000000000000000; // D (0x00000000020000000001000000000000) 
14'h022f : LOC =         127'b0000000000000000000000000000000000001000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000; // D (0x00000000040000000001000000000000) 
14'h2bdb : LOC =         127'b0000000000000000000000000000000000010000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000; // D (0x00000000080000000001000000000000) 
14'h3b44 : LOC =         127'b0000000000000000000000000000000000100000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000; // D (0x00000000100000000001000000000000) 
14'h1a7a : LOC =         127'b0000000000000000000000000000000001000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000; // D (0x00000000200000000001000000000000) 
14'h1b71 : LOC =         127'b0000000000000000000000000000000010000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000; // D (0x00000000400000000001000000000000) 
14'h1967 : LOC =         127'b0000000000000000000000000000000100000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000; // D (0x00000000800000000001000000000000) 
14'h1d4b : LOC =         127'b0000000000000000000000000000001000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000; // D (0x00000001000000000001000000000000) 
14'h1513 : LOC =         127'b0000000000000000000000000000010000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000; // D (0x00000002000000000001000000000000) 
14'h05a3 : LOC =         127'b0000000000000000000000000000100000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000; // D (0x00000004000000000001000000000000) 
14'h24c3 : LOC =         127'b0000000000000000000000000001000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000; // D (0x00000008000000000001000000000000) 
14'h2574 : LOC =         127'b0000000000000000000000000010000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000; // D (0x00000010000000000001000000000000) 
14'h261a : LOC =         127'b0000000000000000000000000100000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000; // D (0x00000020000000000001000000000000) 
14'h20c6 : LOC =         127'b0000000000000000000000001000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000; // D (0x00000040000000000001000000000000) 
14'h2d7e : LOC =         127'b0000000000000000000000010000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000; // D (0x00000080000000000001000000000000) 
14'h360e : LOC =         127'b0000000000000000000000100000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000; // D (0x00000100000000000001000000000000) 
14'h00ee : LOC =         127'b0000000000000000000001000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000; // D (0x00000200000000000001000000000000) 
14'h2e59 : LOC =         127'b0000000000000000000010000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000; // D (0x00000400000000000001000000000000) 
14'h3040 : LOC =         127'b0000000000000000000100000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000; // D (0x00000800000000000001000000000000) 
14'h0c72 : LOC =         127'b0000000000000000001000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000; // D (0x00001000000000000001000000000000) 
14'h3761 : LOC =         127'b0000000000000000010000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000; // D (0x00002000000000000001000000000000) 
14'h0230 : LOC =         127'b0000000000000000100000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000; // D (0x00004000000000000001000000000000) 
14'h2be5 : LOC =         127'b0000000000000001000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000; // D (0x00008000000000000001000000000000) 
14'h3b38 : LOC =         127'b0000000000000010000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000; // D (0x00010000000000000001000000000000) 
14'h1a82 : LOC =         127'b0000000000000100000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000; // D (0x00020000000000000001000000000000) 
14'h1a81 : LOC =         127'b0000000000001000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000; // D (0x00040000000000000001000000000000) 
14'h1a87 : LOC =         127'b0000000000010000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000; // D (0x00080000000000000001000000000000) 
14'h1a8b : LOC =         127'b0000000000100000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000; // D (0x00100000000000000001000000000000) 
14'h1a93 : LOC =         127'b0000000001000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000; // D (0x00200000000000000001000000000000) 
14'h1aa3 : LOC =         127'b0000000010000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000; // D (0x00400000000000000001000000000000) 
14'h1ac3 : LOC =         127'b0000000100000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000; // D (0x00800000000000000001000000000000) 
14'h1a03 : LOC =         127'b0000001000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000; // D (0x01000000000000000001000000000000) 
14'h1b83 : LOC =         127'b0000010000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000; // D (0x02000000000000000001000000000000) 
14'h1883 : LOC =         127'b0000100000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000; // D (0x04000000000000000001000000000000) 
14'h1e83 : LOC =         127'b0001000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000; // D (0x08000000000000000001000000000000) 
14'h1283 : LOC =         127'b0010000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000; // D (0x10000000000000000001000000000000) 
14'h0a83 : LOC =         127'b0100000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000; // D (0x20000000000000000001000000000000) 
14'h3a83 : LOC =         127'b1000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000; // D (0x40000000000000000001000000000000) 
14'h3506 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000; // S (0x00000000000000000002000000000000) 
14'h1c7d : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000000000000000000000000000000; // D (0x00000000000000000006000000000000) 
14'h2487 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000001010000000000000000000000000000000000000000000000000; // D (0x0000000000000000000a000000000000) 
14'h1604 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000; // D (0x00000000000000000012000000000000) 
14'h3075 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000100010000000000000000000000000000000000000000000000000; // D (0x00000000000000000022000000000000) 
14'h3fe0 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000001000010000000000000000000000000000000000000000000000000; // D (0x00000000000000000042000000000000) 
14'h20ca : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000010000010000000000000000000000000000000000000000000000000; // D (0x00000000000000000082000000000000) 
14'h1e9e : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000100000010000000000000000000000000000000000000000000000000; // D (0x00000000000000000102000000000000) 
14'h2141 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000001000000010000000000000000000000000000000000000000000000000; // D (0x00000000000000000202000000000000) 
14'h1d88 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000010000000010000000000000000000000000000000000000000000000000; // D (0x00000000000000000402000000000000) 
14'h276d : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000100000000010000000000000000000000000000000000000000000000000; // D (0x00000000000000000802000000000000) 
14'h11d0 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000001000000000010000000000000000000000000000000000000000000000000; // D (0x00000000000000001002000000000000) 
14'h3fdd : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000010000000000010000000000000000000000000000000000000000000000000; // D (0x00000000000000002002000000000000) 
14'h20b0 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000100000000000010000000000000000000000000000000000000000000000000; // D (0x00000000000000004002000000000000) 
14'h1e6a : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000001000000000000010000000000000000000000000000000000000000000000000; // D (0x00000000000000008002000000000000) 
14'h20a9 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000010000000000000010000000000000000000000000000000000000000000000000; // D (0x00000000000000010002000000000000) 
14'h1e58 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000100000000000000010000000000000000000000000000000000000000000000000; // D (0x00000000000000020002000000000000) 
14'h20cd : LOC =         127'b0000000000000000000000000000000000000000000000000000000000001000000000000000010000000000000000000000000000000000000000000000000; // D (0x00000000000000040002000000000000) 
14'h1e90 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000010000000000000000010000000000000000000000000000000000000000000000000; // D (0x00000000000000080002000000000000) 
14'h215d : LOC =         127'b0000000000000000000000000000000000000000000000000000000000100000000000000000010000000000000000000000000000000000000000000000000; // D (0x00000000000000100002000000000000) 
14'h1db0 : LOC =         127'b0000000000000000000000000000000000000000000000000000000001000000000000000000010000000000000000000000000000000000000000000000000; // D (0x00000000000000200002000000000000) 
14'h271d : LOC =         127'b0000000000000000000000000000000000000000000000000000000010000000000000000000010000000000000000000000000000000000000000000000000; // D (0x00000000000000400002000000000000) 
14'h1130 : LOC =         127'b0000000000000000000000000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000000000000000000; // D (0x00000000000000800002000000000000) 
14'h3e1d : LOC =         127'b0000000000000000000000000000000000000000000000000000001000000000000000000000010000000000000000000000000000000000000000000000000; // D (0x00000000000001000002000000000000) 
14'h2330 : LOC =         127'b0000000000000000000000000000000000000000000000000000010000000000000000000000010000000000000000000000000000000000000000000000000; // D (0x00000000000002000002000000000000) 
14'h196a : LOC =         127'b0000000000000000000000000000000000000000000000000000100000000000000000000000010000000000000000000000000000000000000000000000000; // D (0x00000000000004000002000000000000) 
14'h2ea9 : LOC =         127'b0000000000000000000000000000000000000000000000000001000000000000000000000000010000000000000000000000000000000000000000000000000; // D (0x00000000000008000002000000000000) 
14'h0258 : LOC =         127'b0000000000000000000000000000000000000000000000000010000000000000000000000000010000000000000000000000000000000000000000000000000; // D (0x00000000000010000002000000000000) 
14'h18cd : LOC =         127'b0000000000000000000000000000000000000000000000000100000000000000000000000000010000000000000000000000000000000000000000000000000; // D (0x00000000000020000002000000000000) 
14'h2de7 : LOC =         127'b0000000000000000000000000000000000000000000000001000000000000000000000000000010000000000000000000000000000000000000000000000000; // D (0x00000000000040000002000000000000) 
14'h04c4 : LOC =         127'b0000000000000000000000000000000000000000000000010000000000000000000000000000010000000000000000000000000000000000000000000000000; // D (0x00000000000080000002000000000000) 
14'h15f5 : LOC =         127'b0000000000000000000000000000000000000000000000100000000000000000000000000000010000000000000000000000000000000000000000000000000; // D (0x00000000000100000002000000000000) 
14'h3797 : LOC =         127'b0000000000000000000000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000000000000000000000; // D (0x00000000000200000002000000000000) 
14'h3024 : LOC =         127'b0000000000000000000000000000000000000000000010000000000000000000000000000000010000000000000000000000000000000000000000000000000; // D (0x00000000000400000002000000000000) 
14'h3f42 : LOC =         127'b0000000000000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000000000000000000; // D (0x00000000000800000002000000000000) 
14'h218e : LOC =         127'b0000000000000000000000000000000000000000001000000000000000000000000000000000010000000000000000000000000000000000000000000000000; // D (0x00000000001000000002000000000000) 
14'h1c16 : LOC =         127'b0000000000000000000000000000000000000000010000000000000000000000000000000000010000000000000000000000000000000000000000000000000; // D (0x00000000002000000002000000000000) 
14'h2451 : LOC =         127'b0000000000000000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000000000000000000; // D (0x00000000004000000002000000000000) 
14'h17a8 : LOC =         127'b0000000000000000000000000000000000000001000000000000000000000000000000000000010000000000000000000000000000000000000000000000000; // D (0x00000000008000000002000000000000) 
14'h332d : LOC =         127'b0000000000000000000000000000000000000010000000000000000000000000000000000000010000000000000000000000000000000000000000000000000; // D (0x00000000010000000002000000000000) 
14'h3950 : LOC =         127'b0000000000000000000000000000000000000100000000000000000000000000000000000000010000000000000000000000000000000000000000000000000; // D (0x00000000020000000002000000000000) 
14'h2daa : LOC =         127'b0000000000000000000000000000000000001000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000; // D (0x00000000040000000002000000000000) 
14'h045e : LOC =         127'b0000000000000000000000000000000000010000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000; // D (0x00000000080000000002000000000000) 
14'h14c1 : LOC =         127'b0000000000000000000000000000000000100000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000; // D (0x00000000100000000002000000000000) 
14'h35ff : LOC =         127'b0000000000000000000000000000000001000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000; // D (0x00000000200000000002000000000000) 
14'h34f4 : LOC =         127'b0000000000000000000000000000000010000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000; // D (0x00000000400000000002000000000000) 
14'h36e2 : LOC =         127'b0000000000000000000000000000000100000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000; // D (0x00000000800000000002000000000000) 
14'h32ce : LOC =         127'b0000000000000000000000000000001000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000; // D (0x00000001000000000002000000000000) 
14'h3a96 : LOC =         127'b0000000000000000000000000000010000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000; // D (0x00000002000000000002000000000000) 
14'h2a26 : LOC =         127'b0000000000000000000000000000100000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000; // D (0x00000004000000000002000000000000) 
14'h0b46 : LOC =         127'b0000000000000000000000000001000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000; // D (0x00000008000000000002000000000000) 
14'h0af1 : LOC =         127'b0000000000000000000000000010000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000; // D (0x00000010000000000002000000000000) 
14'h099f : LOC =         127'b0000000000000000000000000100000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000; // D (0x00000020000000000002000000000000) 
14'h0f43 : LOC =         127'b0000000000000000000000001000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000; // D (0x00000040000000000002000000000000) 
14'h02fb : LOC =         127'b0000000000000000000000010000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000; // D (0x00000080000000000002000000000000) 
14'h198b : LOC =         127'b0000000000000000000000100000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000; // D (0x00000100000000000002000000000000) 
14'h2f6b : LOC =         127'b0000000000000000000001000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000; // D (0x00000200000000000002000000000000) 
14'h01dc : LOC =         127'b0000000000000000000010000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000; // D (0x00000400000000000002000000000000) 
14'h1fc5 : LOC =         127'b0000000000000000000100000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000; // D (0x00000800000000000002000000000000) 
14'h23f7 : LOC =         127'b0000000000000000001000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000; // D (0x00001000000000000002000000000000) 
14'h18e4 : LOC =         127'b0000000000000000010000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000; // D (0x00002000000000000002000000000000) 
14'h2db5 : LOC =         127'b0000000000000000100000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000; // D (0x00004000000000000002000000000000) 
14'h0460 : LOC =         127'b0000000000000001000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000; // D (0x00008000000000000002000000000000) 
14'h14bd : LOC =         127'b0000000000000010000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000; // D (0x00010000000000000002000000000000) 
14'h3507 : LOC =         127'b0000000000000100000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000; // D (0x00020000000000000002000000000000) 
14'h3504 : LOC =         127'b0000000000001000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000; // D (0x00040000000000000002000000000000) 
14'h3502 : LOC =         127'b0000000000010000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000; // D (0x00080000000000000002000000000000) 
14'h350e : LOC =         127'b0000000000100000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000; // D (0x00100000000000000002000000000000) 
14'h3516 : LOC =         127'b0000000001000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000; // D (0x00200000000000000002000000000000) 
14'h3526 : LOC =         127'b0000000010000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000; // D (0x00400000000000000002000000000000) 
14'h3546 : LOC =         127'b0000000100000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000; // D (0x00800000000000000002000000000000) 
14'h3586 : LOC =         127'b0000001000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000; // D (0x01000000000000000002000000000000) 
14'h3406 : LOC =         127'b0000010000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000; // D (0x02000000000000000002000000000000) 
14'h3706 : LOC =         127'b0000100000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000; // D (0x04000000000000000002000000000000) 
14'h3106 : LOC =         127'b0001000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000; // D (0x08000000000000000002000000000000) 
14'h3d06 : LOC =         127'b0010000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000; // D (0x10000000000000000002000000000000) 
14'h2506 : LOC =         127'b0100000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000; // D (0x20000000000000000002000000000000) 
14'h1506 : LOC =         127'b1000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000; // D (0x40000000000000000002000000000000) 
14'h297b : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000; // S (0x00000000000000000004000000000000) 
14'h38fa : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000000000000000000000000; // D (0x0000000000000000000c000000000000) 
14'h0a79 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000000000000000000000000000; // D (0x00000000000000000014000000000000) 
14'h2c08 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000; // D (0x00000000000000000024000000000000) 
14'h239d : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000001000100000000000000000000000000000000000000000000000000; // D (0x00000000000000000044000000000000) 
14'h3cb7 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000010000100000000000000000000000000000000000000000000000000; // D (0x00000000000000000084000000000000) 
14'h02e3 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000100000100000000000000000000000000000000000000000000000000; // D (0x00000000000000000104000000000000) 
14'h3d3c : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000001000000100000000000000000000000000000000000000000000000000; // D (0x00000000000000000204000000000000) 
14'h01f5 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000010000000100000000000000000000000000000000000000000000000000; // D (0x00000000000000000404000000000000) 
14'h3b10 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000100000000100000000000000000000000000000000000000000000000000; // D (0x00000000000000000804000000000000) 
14'h0dad : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000001000000000100000000000000000000000000000000000000000000000000; // D (0x00000000000000001004000000000000) 
14'h23a0 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000010000000000100000000000000000000000000000000000000000000000000; // D (0x00000000000000002004000000000000) 
14'h3ccd : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000100000000000100000000000000000000000000000000000000000000000000; // D (0x00000000000000004004000000000000) 
14'h0217 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000001000000000000100000000000000000000000000000000000000000000000000; // D (0x00000000000000008004000000000000) 
14'h3cd4 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000010000000000000100000000000000000000000000000000000000000000000000; // D (0x00000000000000010004000000000000) 
14'h0225 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000100000000000000100000000000000000000000000000000000000000000000000; // D (0x00000000000000020004000000000000) 
14'h3cb0 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000001000000000000000100000000000000000000000000000000000000000000000000; // D (0x00000000000000040004000000000000) 
14'h02ed : LOC =         127'b0000000000000000000000000000000000000000000000000000000000010000000000000000100000000000000000000000000000000000000000000000000; // D (0x00000000000000080004000000000000) 
14'h3d20 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000100000000000000000100000000000000000000000000000000000000000000000000; // D (0x00000000000000100004000000000000) 
14'h01cd : LOC =         127'b0000000000000000000000000000000000000000000000000000000001000000000000000000100000000000000000000000000000000000000000000000000; // D (0x00000000000000200004000000000000) 
14'h3b60 : LOC =         127'b0000000000000000000000000000000000000000000000000000000010000000000000000000100000000000000000000000000000000000000000000000000; // D (0x00000000000000400004000000000000) 
14'h0d4d : LOC =         127'b0000000000000000000000000000000000000000000000000000000100000000000000000000100000000000000000000000000000000000000000000000000; // D (0x00000000000000800004000000000000) 
14'h2260 : LOC =         127'b0000000000000000000000000000000000000000000000000000001000000000000000000000100000000000000000000000000000000000000000000000000; // D (0x00000000000001000004000000000000) 
14'h3f4d : LOC =         127'b0000000000000000000000000000000000000000000000000000010000000000000000000000100000000000000000000000000000000000000000000000000; // D (0x00000000000002000004000000000000) 
14'h0517 : LOC =         127'b0000000000000000000000000000000000000000000000000000100000000000000000000000100000000000000000000000000000000000000000000000000; // D (0x00000000000004000004000000000000) 
14'h32d4 : LOC =         127'b0000000000000000000000000000000000000000000000000001000000000000000000000000100000000000000000000000000000000000000000000000000; // D (0x00000000000008000004000000000000) 
14'h1e25 : LOC =         127'b0000000000000000000000000000000000000000000000000010000000000000000000000000100000000000000000000000000000000000000000000000000; // D (0x00000000000010000004000000000000) 
14'h04b0 : LOC =         127'b0000000000000000000000000000000000000000000000000100000000000000000000000000100000000000000000000000000000000000000000000000000; // D (0x00000000000020000004000000000000) 
14'h319a : LOC =         127'b0000000000000000000000000000000000000000000000001000000000000000000000000000100000000000000000000000000000000000000000000000000; // D (0x00000000000040000004000000000000) 
14'h18b9 : LOC =         127'b0000000000000000000000000000000000000000000000010000000000000000000000000000100000000000000000000000000000000000000000000000000; // D (0x00000000000080000004000000000000) 
14'h0988 : LOC =         127'b0000000000000000000000000000000000000000000000100000000000000000000000000000100000000000000000000000000000000000000000000000000; // D (0x00000000000100000004000000000000) 
14'h2bea : LOC =         127'b0000000000000000000000000000000000000000000001000000000000000000000000000000100000000000000000000000000000000000000000000000000; // D (0x00000000000200000004000000000000) 
14'h2c59 : LOC =         127'b0000000000000000000000000000000000000000000010000000000000000000000000000000100000000000000000000000000000000000000000000000000; // D (0x00000000000400000004000000000000) 
14'h233f : LOC =         127'b0000000000000000000000000000000000000000000100000000000000000000000000000000100000000000000000000000000000000000000000000000000; // D (0x00000000000800000004000000000000) 
14'h3df3 : LOC =         127'b0000000000000000000000000000000000000000001000000000000000000000000000000000100000000000000000000000000000000000000000000000000; // D (0x00000000001000000004000000000000) 
14'h006b : LOC =         127'b0000000000000000000000000000000000000000010000000000000000000000000000000000100000000000000000000000000000000000000000000000000; // D (0x00000000002000000004000000000000) 
14'h382c : LOC =         127'b0000000000000000000000000000000000000000100000000000000000000000000000000000100000000000000000000000000000000000000000000000000; // D (0x00000000004000000004000000000000) 
14'h0bd5 : LOC =         127'b0000000000000000000000000000000000000001000000000000000000000000000000000000100000000000000000000000000000000000000000000000000; // D (0x00000000008000000004000000000000) 
14'h2f50 : LOC =         127'b0000000000000000000000000000000000000010000000000000000000000000000000000000100000000000000000000000000000000000000000000000000; // D (0x00000000010000000004000000000000) 
14'h252d : LOC =         127'b0000000000000000000000000000000000000100000000000000000000000000000000000000100000000000000000000000000000000000000000000000000; // D (0x00000000020000000004000000000000) 
14'h31d7 : LOC =         127'b0000000000000000000000000000000000001000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000; // D (0x00000000040000000004000000000000) 
14'h1823 : LOC =         127'b0000000000000000000000000000000000010000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000; // D (0x00000000080000000004000000000000) 
14'h08bc : LOC =         127'b0000000000000000000000000000000000100000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000; // D (0x00000000100000000004000000000000) 
14'h2982 : LOC =         127'b0000000000000000000000000000000001000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000; // D (0x00000000200000000004000000000000) 
14'h2889 : LOC =         127'b0000000000000000000000000000000010000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000; // D (0x00000000400000000004000000000000) 
14'h2a9f : LOC =         127'b0000000000000000000000000000000100000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000; // D (0x00000000800000000004000000000000) 
14'h2eb3 : LOC =         127'b0000000000000000000000000000001000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000; // D (0x00000001000000000004000000000000) 
14'h26eb : LOC =         127'b0000000000000000000000000000010000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000; // D (0x00000002000000000004000000000000) 
14'h365b : LOC =         127'b0000000000000000000000000000100000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000; // D (0x00000004000000000004000000000000) 
14'h173b : LOC =         127'b0000000000000000000000000001000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000; // D (0x00000008000000000004000000000000) 
14'h168c : LOC =         127'b0000000000000000000000000010000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000; // D (0x00000010000000000004000000000000) 
14'h15e2 : LOC =         127'b0000000000000000000000000100000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000; // D (0x00000020000000000004000000000000) 
14'h133e : LOC =         127'b0000000000000000000000001000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000; // D (0x00000040000000000004000000000000) 
14'h1e86 : LOC =         127'b0000000000000000000000010000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000; // D (0x00000080000000000004000000000000) 
14'h05f6 : LOC =         127'b0000000000000000000000100000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000; // D (0x00000100000000000004000000000000) 
14'h3316 : LOC =         127'b0000000000000000000001000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000; // D (0x00000200000000000004000000000000) 
14'h1da1 : LOC =         127'b0000000000000000000010000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000; // D (0x00000400000000000004000000000000) 
14'h03b8 : LOC =         127'b0000000000000000000100000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000; // D (0x00000800000000000004000000000000) 
14'h3f8a : LOC =         127'b0000000000000000001000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000; // D (0x00001000000000000004000000000000) 
14'h0499 : LOC =         127'b0000000000000000010000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000; // D (0x00002000000000000004000000000000) 
14'h31c8 : LOC =         127'b0000000000000000100000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000; // D (0x00004000000000000004000000000000) 
14'h181d : LOC =         127'b0000000000000001000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000; // D (0x00008000000000000004000000000000) 
14'h08c0 : LOC =         127'b0000000000000010000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000; // D (0x00010000000000000004000000000000) 
14'h297a : LOC =         127'b0000000000000100000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000; // D (0x00020000000000000004000000000000) 
14'h2979 : LOC =         127'b0000000000001000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000; // D (0x00040000000000000004000000000000) 
14'h297f : LOC =         127'b0000000000010000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000; // D (0x00080000000000000004000000000000) 
14'h2973 : LOC =         127'b0000000000100000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000; // D (0x00100000000000000004000000000000) 
14'h296b : LOC =         127'b0000000001000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000; // D (0x00200000000000000004000000000000) 
14'h295b : LOC =         127'b0000000010000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000; // D (0x00400000000000000004000000000000) 
14'h293b : LOC =         127'b0000000100000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000; // D (0x00800000000000000004000000000000) 
14'h29fb : LOC =         127'b0000001000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000; // D (0x01000000000000000004000000000000) 
14'h287b : LOC =         127'b0000010000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000; // D (0x02000000000000000004000000000000) 
14'h2b7b : LOC =         127'b0000100000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000; // D (0x04000000000000000004000000000000) 
14'h2d7b : LOC =         127'b0001000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000; // D (0x08000000000000000004000000000000) 
14'h217b : LOC =         127'b0010000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000; // D (0x10000000000000000004000000000000) 
14'h397b : LOC =         127'b0100000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000; // D (0x20000000000000000004000000000000) 
14'h097b : LOC =         127'b1000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000; // D (0x40000000000000000004000000000000) 
14'h1181 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000; // S (0x00000000000000000008000000000000) 
14'h3283 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000000000000000000000000000000; // D (0x00000000000000000018000000000000) 
14'h14f2 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000101000000000000000000000000000000000000000000000000000; // D (0x00000000000000000028000000000000) 
14'h1b67 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000; // D (0x00000000000000000048000000000000) 
14'h044d : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000010001000000000000000000000000000000000000000000000000000; // D (0x00000000000000000088000000000000) 
14'h3a19 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000100001000000000000000000000000000000000000000000000000000; // D (0x00000000000000000108000000000000) 
14'h05c6 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000001000001000000000000000000000000000000000000000000000000000; // D (0x00000000000000000208000000000000) 
14'h390f : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000010000001000000000000000000000000000000000000000000000000000; // D (0x00000000000000000408000000000000) 
14'h03ea : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000100000001000000000000000000000000000000000000000000000000000; // D (0x00000000000000000808000000000000) 
14'h3557 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000001000000001000000000000000000000000000000000000000000000000000; // D (0x00000000000000001008000000000000) 
14'h1b5a : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000010000000001000000000000000000000000000000000000000000000000000; // D (0x00000000000000002008000000000000) 
14'h0437 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000100000000001000000000000000000000000000000000000000000000000000; // D (0x00000000000000004008000000000000) 
14'h3aed : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000001000000000001000000000000000000000000000000000000000000000000000; // D (0x00000000000000008008000000000000) 
14'h042e : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000010000000000001000000000000000000000000000000000000000000000000000; // D (0x00000000000000010008000000000000) 
14'h3adf : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000100000000000001000000000000000000000000000000000000000000000000000; // D (0x00000000000000020008000000000000) 
14'h044a : LOC =         127'b0000000000000000000000000000000000000000000000000000000000001000000000000001000000000000000000000000000000000000000000000000000; // D (0x00000000000000040008000000000000) 
14'h3a17 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000010000000000000001000000000000000000000000000000000000000000000000000; // D (0x00000000000000080008000000000000) 
14'h05da : LOC =         127'b0000000000000000000000000000000000000000000000000000000000100000000000000001000000000000000000000000000000000000000000000000000; // D (0x00000000000000100008000000000000) 
14'h3937 : LOC =         127'b0000000000000000000000000000000000000000000000000000000001000000000000000001000000000000000000000000000000000000000000000000000; // D (0x00000000000000200008000000000000) 
14'h039a : LOC =         127'b0000000000000000000000000000000000000000000000000000000010000000000000000001000000000000000000000000000000000000000000000000000; // D (0x00000000000000400008000000000000) 
14'h35b7 : LOC =         127'b0000000000000000000000000000000000000000000000000000000100000000000000000001000000000000000000000000000000000000000000000000000; // D (0x00000000000000800008000000000000) 
14'h1a9a : LOC =         127'b0000000000000000000000000000000000000000000000000000001000000000000000000001000000000000000000000000000000000000000000000000000; // D (0x00000000000001000008000000000000) 
14'h07b7 : LOC =         127'b0000000000000000000000000000000000000000000000000000010000000000000000000001000000000000000000000000000000000000000000000000000; // D (0x00000000000002000008000000000000) 
14'h3ded : LOC =         127'b0000000000000000000000000000000000000000000000000000100000000000000000000001000000000000000000000000000000000000000000000000000; // D (0x00000000000004000008000000000000) 
14'h0a2e : LOC =         127'b0000000000000000000000000000000000000000000000000001000000000000000000000001000000000000000000000000000000000000000000000000000; // D (0x00000000000008000008000000000000) 
14'h26df : LOC =         127'b0000000000000000000000000000000000000000000000000010000000000000000000000001000000000000000000000000000000000000000000000000000; // D (0x00000000000010000008000000000000) 
14'h3c4a : LOC =         127'b0000000000000000000000000000000000000000000000000100000000000000000000000001000000000000000000000000000000000000000000000000000; // D (0x00000000000020000008000000000000) 
14'h0960 : LOC =         127'b0000000000000000000000000000000000000000000000001000000000000000000000000001000000000000000000000000000000000000000000000000000; // D (0x00000000000040000008000000000000) 
14'h2043 : LOC =         127'b0000000000000000000000000000000000000000000000010000000000000000000000000001000000000000000000000000000000000000000000000000000; // D (0x00000000000080000008000000000000) 
14'h3172 : LOC =         127'b0000000000000000000000000000000000000000000000100000000000000000000000000001000000000000000000000000000000000000000000000000000; // D (0x00000000000100000008000000000000) 
14'h1310 : LOC =         127'b0000000000000000000000000000000000000000000001000000000000000000000000000001000000000000000000000000000000000000000000000000000; // D (0x00000000000200000008000000000000) 
14'h14a3 : LOC =         127'b0000000000000000000000000000000000000000000010000000000000000000000000000001000000000000000000000000000000000000000000000000000; // D (0x00000000000400000008000000000000) 
14'h1bc5 : LOC =         127'b0000000000000000000000000000000000000000000100000000000000000000000000000001000000000000000000000000000000000000000000000000000; // D (0x00000000000800000008000000000000) 
14'h0509 : LOC =         127'b0000000000000000000000000000000000000000001000000000000000000000000000000001000000000000000000000000000000000000000000000000000; // D (0x00000000001000000008000000000000) 
14'h3891 : LOC =         127'b0000000000000000000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000000000000000000000000; // D (0x00000000002000000008000000000000) 
14'h00d6 : LOC =         127'b0000000000000000000000000000000000000000100000000000000000000000000000000001000000000000000000000000000000000000000000000000000; // D (0x00000000004000000008000000000000) 
14'h332f : LOC =         127'b0000000000000000000000000000000000000001000000000000000000000000000000000001000000000000000000000000000000000000000000000000000; // D (0x00000000008000000008000000000000) 
14'h17aa : LOC =         127'b0000000000000000000000000000000000000010000000000000000000000000000000000001000000000000000000000000000000000000000000000000000; // D (0x00000000010000000008000000000000) 
14'h1dd7 : LOC =         127'b0000000000000000000000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000000000000000000; // D (0x00000000020000000008000000000000) 
14'h092d : LOC =         127'b0000000000000000000000000000000000001000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000; // D (0x00000000040000000008000000000000) 
14'h20d9 : LOC =         127'b0000000000000000000000000000000000010000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000; // D (0x00000000080000000008000000000000) 
14'h3046 : LOC =         127'b0000000000000000000000000000000000100000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000; // D (0x00000000100000000008000000000000) 
14'h1178 : LOC =         127'b0000000000000000000000000000000001000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000; // D (0x00000000200000000008000000000000) 
14'h1073 : LOC =         127'b0000000000000000000000000000000010000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000; // D (0x00000000400000000008000000000000) 
14'h1265 : LOC =         127'b0000000000000000000000000000000100000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000; // D (0x00000000800000000008000000000000) 
14'h1649 : LOC =         127'b0000000000000000000000000000001000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000; // D (0x00000001000000000008000000000000) 
14'h1e11 : LOC =         127'b0000000000000000000000000000010000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000; // D (0x00000002000000000008000000000000) 
14'h0ea1 : LOC =         127'b0000000000000000000000000000100000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000; // D (0x00000004000000000008000000000000) 
14'h2fc1 : LOC =         127'b0000000000000000000000000001000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000; // D (0x00000008000000000008000000000000) 
14'h2e76 : LOC =         127'b0000000000000000000000000010000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000; // D (0x00000010000000000008000000000000) 
14'h2d18 : LOC =         127'b0000000000000000000000000100000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000; // D (0x00000020000000000008000000000000) 
14'h2bc4 : LOC =         127'b0000000000000000000000001000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000; // D (0x00000040000000000008000000000000) 
14'h267c : LOC =         127'b0000000000000000000000010000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000; // D (0x00000080000000000008000000000000) 
14'h3d0c : LOC =         127'b0000000000000000000000100000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000; // D (0x00000100000000000008000000000000) 
14'h0bec : LOC =         127'b0000000000000000000001000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000; // D (0x00000200000000000008000000000000) 
14'h255b : LOC =         127'b0000000000000000000010000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000; // D (0x00000400000000000008000000000000) 
14'h3b42 : LOC =         127'b0000000000000000000100000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000; // D (0x00000800000000000008000000000000) 
14'h0770 : LOC =         127'b0000000000000000001000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000; // D (0x00001000000000000008000000000000) 
14'h3c63 : LOC =         127'b0000000000000000010000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000; // D (0x00002000000000000008000000000000) 
14'h0932 : LOC =         127'b0000000000000000100000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000; // D (0x00004000000000000008000000000000) 
14'h20e7 : LOC =         127'b0000000000000001000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000; // D (0x00008000000000000008000000000000) 
14'h303a : LOC =         127'b0000000000000010000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000; // D (0x00010000000000000008000000000000) 
14'h1180 : LOC =         127'b0000000000000100000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000; // D (0x00020000000000000008000000000000) 
14'h1183 : LOC =         127'b0000000000001000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000; // D (0x00040000000000000008000000000000) 
14'h1185 : LOC =         127'b0000000000010000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000; // D (0x00080000000000000008000000000000) 
14'h1189 : LOC =         127'b0000000000100000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000; // D (0x00100000000000000008000000000000) 
14'h1191 : LOC =         127'b0000000001000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000; // D (0x00200000000000000008000000000000) 
14'h11a1 : LOC =         127'b0000000010000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000; // D (0x00400000000000000008000000000000) 
14'h11c1 : LOC =         127'b0000000100000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000; // D (0x00800000000000000008000000000000) 
14'h1101 : LOC =         127'b0000001000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000; // D (0x01000000000000000008000000000000) 
14'h1081 : LOC =         127'b0000010000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000; // D (0x02000000000000000008000000000000) 
14'h1381 : LOC =         127'b0000100000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000; // D (0x04000000000000000008000000000000) 
14'h1581 : LOC =         127'b0001000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000; // D (0x08000000000000000008000000000000) 
14'h1981 : LOC =         127'b0010000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000; // D (0x10000000000000000008000000000000) 
14'h0181 : LOC =         127'b0100000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000; // D (0x20000000000000000008000000000000) 
14'h3181 : LOC =         127'b1000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000; // D (0x40000000000000000008000000000000) 
14'h2302 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000; // S (0x00000000000000000010000000000000) 
14'h2671 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000000000000000000000000000000000; // D (0x00000000000000000030000000000000) 
14'h29e4 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000001010000000000000000000000000000000000000000000000000000; // D (0x00000000000000000050000000000000) 
14'h36ce : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000; // D (0x00000000000000000090000000000000) 
14'h089a : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000100010000000000000000000000000000000000000000000000000000; // D (0x00000000000000000110000000000000) 
14'h3745 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000001000010000000000000000000000000000000000000000000000000000; // D (0x00000000000000000210000000000000) 
14'h0b8c : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000010000010000000000000000000000000000000000000000000000000000; // D (0x00000000000000000410000000000000) 
14'h3169 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000100000010000000000000000000000000000000000000000000000000000; // D (0x00000000000000000810000000000000) 
14'h07d4 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000001000000010000000000000000000000000000000000000000000000000000; // D (0x00000000000000001010000000000000) 
14'h29d9 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000010000000010000000000000000000000000000000000000000000000000000; // D (0x00000000000000002010000000000000) 
14'h36b4 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000100000000010000000000000000000000000000000000000000000000000000; // D (0x00000000000000004010000000000000) 
14'h086e : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000001000000000010000000000000000000000000000000000000000000000000000; // D (0x00000000000000008010000000000000) 
14'h36ad : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000010000000000010000000000000000000000000000000000000000000000000000; // D (0x00000000000000010010000000000000) 
14'h085c : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000100000000000010000000000000000000000000000000000000000000000000000; // D (0x00000000000000020010000000000000) 
14'h36c9 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000001000000000000010000000000000000000000000000000000000000000000000000; // D (0x00000000000000040010000000000000) 
14'h0894 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000010000000000000010000000000000000000000000000000000000000000000000000; // D (0x00000000000000080010000000000000) 
14'h3759 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000100000000000000010000000000000000000000000000000000000000000000000000; // D (0x00000000000000100010000000000000) 
14'h0bb4 : LOC =         127'b0000000000000000000000000000000000000000000000000000000001000000000000000010000000000000000000000000000000000000000000000000000; // D (0x00000000000000200010000000000000) 
14'h3119 : LOC =         127'b0000000000000000000000000000000000000000000000000000000010000000000000000010000000000000000000000000000000000000000000000000000; // D (0x00000000000000400010000000000000) 
14'h0734 : LOC =         127'b0000000000000000000000000000000000000000000000000000000100000000000000000010000000000000000000000000000000000000000000000000000; // D (0x00000000000000800010000000000000) 
14'h2819 : LOC =         127'b0000000000000000000000000000000000000000000000000000001000000000000000000010000000000000000000000000000000000000000000000000000; // D (0x00000000000001000010000000000000) 
14'h3534 : LOC =         127'b0000000000000000000000000000000000000000000000000000010000000000000000000010000000000000000000000000000000000000000000000000000; // D (0x00000000000002000010000000000000) 
14'h0f6e : LOC =         127'b0000000000000000000000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000000000000000000000; // D (0x00000000000004000010000000000000) 
14'h38ad : LOC =         127'b0000000000000000000000000000000000000000000000000001000000000000000000000010000000000000000000000000000000000000000000000000000; // D (0x00000000000008000010000000000000) 
14'h145c : LOC =         127'b0000000000000000000000000000000000000000000000000010000000000000000000000010000000000000000000000000000000000000000000000000000; // D (0x00000000000010000010000000000000) 
14'h0ec9 : LOC =         127'b0000000000000000000000000000000000000000000000000100000000000000000000000010000000000000000000000000000000000000000000000000000; // D (0x00000000000020000010000000000000) 
14'h3be3 : LOC =         127'b0000000000000000000000000000000000000000000000001000000000000000000000000010000000000000000000000000000000000000000000000000000; // D (0x00000000000040000010000000000000) 
14'h12c0 : LOC =         127'b0000000000000000000000000000000000000000000000010000000000000000000000000010000000000000000000000000000000000000000000000000000; // D (0x00000000000080000010000000000000) 
14'h03f1 : LOC =         127'b0000000000000000000000000000000000000000000000100000000000000000000000000010000000000000000000000000000000000000000000000000000; // D (0x00000000000100000010000000000000) 
14'h2193 : LOC =         127'b0000000000000000000000000000000000000000000001000000000000000000000000000010000000000000000000000000000000000000000000000000000; // D (0x00000000000200000010000000000000) 
14'h2620 : LOC =         127'b0000000000000000000000000000000000000000000010000000000000000000000000000010000000000000000000000000000000000000000000000000000; // D (0x00000000000400000010000000000000) 
14'h2946 : LOC =         127'b0000000000000000000000000000000000000000000100000000000000000000000000000010000000000000000000000000000000000000000000000000000; // D (0x00000000000800000010000000000000) 
14'h378a : LOC =         127'b0000000000000000000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000000000000000000000000; // D (0x00000000001000000010000000000000) 
14'h0a12 : LOC =         127'b0000000000000000000000000000000000000000010000000000000000000000000000000010000000000000000000000000000000000000000000000000000; // D (0x00000000002000000010000000000000) 
14'h3255 : LOC =         127'b0000000000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000000000000000000000; // D (0x00000000004000000010000000000000) 
14'h01ac : LOC =         127'b0000000000000000000000000000000000000001000000000000000000000000000000000010000000000000000000000000000000000000000000000000000; // D (0x00000000008000000010000000000000) 
14'h2529 : LOC =         127'b0000000000000000000000000000000000000010000000000000000000000000000000000010000000000000000000000000000000000000000000000000000; // D (0x00000000010000000010000000000000) 
14'h2f54 : LOC =         127'b0000000000000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000000000000000000000; // D (0x00000000020000000010000000000000) 
14'h3bae : LOC =         127'b0000000000000000000000000000000000001000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000; // D (0x00000000040000000010000000000000) 
14'h125a : LOC =         127'b0000000000000000000000000000000000010000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000; // D (0x00000000080000000010000000000000) 
14'h02c5 : LOC =         127'b0000000000000000000000000000000000100000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000; // D (0x00000000100000000010000000000000) 
14'h23fb : LOC =         127'b0000000000000000000000000000000001000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000; // D (0x00000000200000000010000000000000) 
14'h22f0 : LOC =         127'b0000000000000000000000000000000010000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000; // D (0x00000000400000000010000000000000) 
14'h20e6 : LOC =         127'b0000000000000000000000000000000100000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000; // D (0x00000000800000000010000000000000) 
14'h24ca : LOC =         127'b0000000000000000000000000000001000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000; // D (0x00000001000000000010000000000000) 
14'h2c92 : LOC =         127'b0000000000000000000000000000010000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000; // D (0x00000002000000000010000000000000) 
14'h3c22 : LOC =         127'b0000000000000000000000000000100000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000; // D (0x00000004000000000010000000000000) 
14'h1d42 : LOC =         127'b0000000000000000000000000001000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000; // D (0x00000008000000000010000000000000) 
14'h1cf5 : LOC =         127'b0000000000000000000000000010000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000; // D (0x00000010000000000010000000000000) 
14'h1f9b : LOC =         127'b0000000000000000000000000100000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000; // D (0x00000020000000000010000000000000) 
14'h1947 : LOC =         127'b0000000000000000000000001000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000; // D (0x00000040000000000010000000000000) 
14'h14ff : LOC =         127'b0000000000000000000000010000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000; // D (0x00000080000000000010000000000000) 
14'h0f8f : LOC =         127'b0000000000000000000000100000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000; // D (0x00000100000000000010000000000000) 
14'h396f : LOC =         127'b0000000000000000000001000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000; // D (0x00000200000000000010000000000000) 
14'h17d8 : LOC =         127'b0000000000000000000010000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000; // D (0x00000400000000000010000000000000) 
14'h09c1 : LOC =         127'b0000000000000000000100000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000; // D (0x00000800000000000010000000000000) 
14'h35f3 : LOC =         127'b0000000000000000001000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000; // D (0x00001000000000000010000000000000) 
14'h0ee0 : LOC =         127'b0000000000000000010000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000; // D (0x00002000000000000010000000000000) 
14'h3bb1 : LOC =         127'b0000000000000000100000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000; // D (0x00004000000000000010000000000000) 
14'h1264 : LOC =         127'b0000000000000001000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000; // D (0x00008000000000000010000000000000) 
14'h02b9 : LOC =         127'b0000000000000010000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000; // D (0x00010000000000000010000000000000) 
14'h2303 : LOC =         127'b0000000000000100000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000; // D (0x00020000000000000010000000000000) 
14'h2300 : LOC =         127'b0000000000001000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000; // D (0x00040000000000000010000000000000) 
14'h2306 : LOC =         127'b0000000000010000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000; // D (0x00080000000000000010000000000000) 
14'h230a : LOC =         127'b0000000000100000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000; // D (0x00100000000000000010000000000000) 
14'h2312 : LOC =         127'b0000000001000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000; // D (0x00200000000000000010000000000000) 
14'h2322 : LOC =         127'b0000000010000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000; // D (0x00400000000000000010000000000000) 
14'h2342 : LOC =         127'b0000000100000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000; // D (0x00800000000000000010000000000000) 
14'h2382 : LOC =         127'b0000001000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000; // D (0x01000000000000000010000000000000) 
14'h2202 : LOC =         127'b0000010000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000; // D (0x02000000000000000010000000000000) 
14'h2102 : LOC =         127'b0000100000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000; // D (0x04000000000000000010000000000000) 
14'h2702 : LOC =         127'b0001000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000; // D (0x08000000000000000010000000000000) 
14'h2b02 : LOC =         127'b0010000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000; // D (0x10000000000000000010000000000000) 
14'h3302 : LOC =         127'b0100000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000; // D (0x20000000000000000010000000000000) 
14'h0302 : LOC =         127'b1000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000; // D (0x40000000000000000010000000000000) 
14'h0573 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000; // S (0x00000000000000000020000000000000) 
14'h0f95 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000; // D (0x00000000000000000060000000000000) 
14'h10bf : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000000000000000000000000000000; // D (0x000000000000000000a0000000000000) 
14'h2eeb : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000; // D (0x00000000000000000120000000000000) 
14'h1134 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000001000100000000000000000000000000000000000000000000000000000; // D (0x00000000000000000220000000000000) 
14'h2dfd : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000010000100000000000000000000000000000000000000000000000000000; // D (0x00000000000000000420000000000000) 
14'h1718 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000100000100000000000000000000000000000000000000000000000000000; // D (0x00000000000000000820000000000000) 
14'h21a5 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000001000000100000000000000000000000000000000000000000000000000000; // D (0x00000000000000001020000000000000) 
14'h0fa8 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000010000000100000000000000000000000000000000000000000000000000000; // D (0x00000000000000002020000000000000) 
14'h10c5 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000100000000100000000000000000000000000000000000000000000000000000; // D (0x00000000000000004020000000000000) 
14'h2e1f : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000001000000000100000000000000000000000000000000000000000000000000000; // D (0x00000000000000008020000000000000) 
14'h10dc : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000010000000000100000000000000000000000000000000000000000000000000000; // D (0x00000000000000010020000000000000) 
14'h2e2d : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000100000000000100000000000000000000000000000000000000000000000000000; // D (0x00000000000000020020000000000000) 
14'h10b8 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000001000000000000100000000000000000000000000000000000000000000000000000; // D (0x00000000000000040020000000000000) 
14'h2ee5 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000010000000000000100000000000000000000000000000000000000000000000000000; // D (0x00000000000000080020000000000000) 
14'h1128 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000100000000000000100000000000000000000000000000000000000000000000000000; // D (0x00000000000000100020000000000000) 
14'h2dc5 : LOC =         127'b0000000000000000000000000000000000000000000000000000000001000000000000000100000000000000000000000000000000000000000000000000000; // D (0x00000000000000200020000000000000) 
14'h1768 : LOC =         127'b0000000000000000000000000000000000000000000000000000000010000000000000000100000000000000000000000000000000000000000000000000000; // D (0x00000000000000400020000000000000) 
14'h2145 : LOC =         127'b0000000000000000000000000000000000000000000000000000000100000000000000000100000000000000000000000000000000000000000000000000000; // D (0x00000000000000800020000000000000) 
14'h0e68 : LOC =         127'b0000000000000000000000000000000000000000000000000000001000000000000000000100000000000000000000000000000000000000000000000000000; // D (0x00000000000001000020000000000000) 
14'h1345 : LOC =         127'b0000000000000000000000000000000000000000000000000000010000000000000000000100000000000000000000000000000000000000000000000000000; // D (0x00000000000002000020000000000000) 
14'h291f : LOC =         127'b0000000000000000000000000000000000000000000000000000100000000000000000000100000000000000000000000000000000000000000000000000000; // D (0x00000000000004000020000000000000) 
14'h1edc : LOC =         127'b0000000000000000000000000000000000000000000000000001000000000000000000000100000000000000000000000000000000000000000000000000000; // D (0x00000000000008000020000000000000) 
14'h322d : LOC =         127'b0000000000000000000000000000000000000000000000000010000000000000000000000100000000000000000000000000000000000000000000000000000; // D (0x00000000000010000020000000000000) 
14'h28b8 : LOC =         127'b0000000000000000000000000000000000000000000000000100000000000000000000000100000000000000000000000000000000000000000000000000000; // D (0x00000000000020000020000000000000) 
14'h1d92 : LOC =         127'b0000000000000000000000000000000000000000000000001000000000000000000000000100000000000000000000000000000000000000000000000000000; // D (0x00000000000040000020000000000000) 
14'h34b1 : LOC =         127'b0000000000000000000000000000000000000000000000010000000000000000000000000100000000000000000000000000000000000000000000000000000; // D (0x00000000000080000020000000000000) 
14'h2580 : LOC =         127'b0000000000000000000000000000000000000000000000100000000000000000000000000100000000000000000000000000000000000000000000000000000; // D (0x00000000000100000020000000000000) 
14'h07e2 : LOC =         127'b0000000000000000000000000000000000000000000001000000000000000000000000000100000000000000000000000000000000000000000000000000000; // D (0x00000000000200000020000000000000) 
14'h0051 : LOC =         127'b0000000000000000000000000000000000000000000010000000000000000000000000000100000000000000000000000000000000000000000000000000000; // D (0x00000000000400000020000000000000) 
14'h0f37 : LOC =         127'b0000000000000000000000000000000000000000000100000000000000000000000000000100000000000000000000000000000000000000000000000000000; // D (0x00000000000800000020000000000000) 
14'h11fb : LOC =         127'b0000000000000000000000000000000000000000001000000000000000000000000000000100000000000000000000000000000000000000000000000000000; // D (0x00000000001000000020000000000000) 
14'h2c63 : LOC =         127'b0000000000000000000000000000000000000000010000000000000000000000000000000100000000000000000000000000000000000000000000000000000; // D (0x00000000002000000020000000000000) 
14'h1424 : LOC =         127'b0000000000000000000000000000000000000000100000000000000000000000000000000100000000000000000000000000000000000000000000000000000; // D (0x00000000004000000020000000000000) 
14'h27dd : LOC =         127'b0000000000000000000000000000000000000001000000000000000000000000000000000100000000000000000000000000000000000000000000000000000; // D (0x00000000008000000020000000000000) 
14'h0358 : LOC =         127'b0000000000000000000000000000000000000010000000000000000000000000000000000100000000000000000000000000000000000000000000000000000; // D (0x00000000010000000020000000000000) 
14'h0925 : LOC =         127'b0000000000000000000000000000000000000100000000000000000000000000000000000100000000000000000000000000000000000000000000000000000; // D (0x00000000020000000020000000000000) 
14'h1ddf : LOC =         127'b0000000000000000000000000000000000001000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000; // D (0x00000000040000000020000000000000) 
14'h342b : LOC =         127'b0000000000000000000000000000000000010000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000; // D (0x00000000080000000020000000000000) 
14'h24b4 : LOC =         127'b0000000000000000000000000000000000100000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000; // D (0x00000000100000000020000000000000) 
14'h058a : LOC =         127'b0000000000000000000000000000000001000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000; // D (0x00000000200000000020000000000000) 
14'h0481 : LOC =         127'b0000000000000000000000000000000010000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000; // D (0x00000000400000000020000000000000) 
14'h0697 : LOC =         127'b0000000000000000000000000000000100000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000; // D (0x00000000800000000020000000000000) 
14'h02bb : LOC =         127'b0000000000000000000000000000001000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000; // D (0x00000001000000000020000000000000) 
14'h0ae3 : LOC =         127'b0000000000000000000000000000010000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000; // D (0x00000002000000000020000000000000) 
14'h1a53 : LOC =         127'b0000000000000000000000000000100000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000; // D (0x00000004000000000020000000000000) 
14'h3b33 : LOC =         127'b0000000000000000000000000001000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000; // D (0x00000008000000000020000000000000) 
14'h3a84 : LOC =         127'b0000000000000000000000000010000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000; // D (0x00000010000000000020000000000000) 
14'h39ea : LOC =         127'b0000000000000000000000000100000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000; // D (0x00000020000000000020000000000000) 
14'h3f36 : LOC =         127'b0000000000000000000000001000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000; // D (0x00000040000000000020000000000000) 
14'h328e : LOC =         127'b0000000000000000000000010000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000; // D (0x00000080000000000020000000000000) 
14'h29fe : LOC =         127'b0000000000000000000000100000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000; // D (0x00000100000000000020000000000000) 
14'h1f1e : LOC =         127'b0000000000000000000001000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000; // D (0x00000200000000000020000000000000) 
14'h31a9 : LOC =         127'b0000000000000000000010000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000; // D (0x00000400000000000020000000000000) 
14'h2fb0 : LOC =         127'b0000000000000000000100000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000; // D (0x00000800000000000020000000000000) 
14'h1382 : LOC =         127'b0000000000000000001000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000; // D (0x00001000000000000020000000000000) 
14'h2891 : LOC =         127'b0000000000000000010000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000; // D (0x00002000000000000020000000000000) 
14'h1dc0 : LOC =         127'b0000000000000000100000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000; // D (0x00004000000000000020000000000000) 
14'h3415 : LOC =         127'b0000000000000001000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000; // D (0x00008000000000000020000000000000) 
14'h24c8 : LOC =         127'b0000000000000010000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000; // D (0x00010000000000000020000000000000) 
14'h0572 : LOC =         127'b0000000000000100000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000; // D (0x00020000000000000020000000000000) 
14'h0571 : LOC =         127'b0000000000001000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000; // D (0x00040000000000000020000000000000) 
14'h0577 : LOC =         127'b0000000000010000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000; // D (0x00080000000000000020000000000000) 
14'h057b : LOC =         127'b0000000000100000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000; // D (0x00100000000000000020000000000000) 
14'h0563 : LOC =         127'b0000000001000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000; // D (0x00200000000000000020000000000000) 
14'h0553 : LOC =         127'b0000000010000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000; // D (0x00400000000000000020000000000000) 
14'h0533 : LOC =         127'b0000000100000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000; // D (0x00800000000000000020000000000000) 
14'h05f3 : LOC =         127'b0000001000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000; // D (0x01000000000000000020000000000000) 
14'h0473 : LOC =         127'b0000010000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000; // D (0x02000000000000000020000000000000) 
14'h0773 : LOC =         127'b0000100000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000; // D (0x04000000000000000020000000000000) 
14'h0173 : LOC =         127'b0001000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000; // D (0x08000000000000000020000000000000) 
14'h0d73 : LOC =         127'b0010000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000; // D (0x10000000000000000020000000000000) 
14'h1573 : LOC =         127'b0100000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000; // D (0x20000000000000000020000000000000) 
14'h2573 : LOC =         127'b1000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000; // D (0x40000000000000000020000000000000) 
14'h0ae6 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000; // S (0x00000000000000000040000000000000) 
14'h1f2a : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000000000000000000000000000000000; // D (0x000000000000000000c0000000000000) 
14'h217e : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000101000000000000000000000000000000000000000000000000000000; // D (0x00000000000000000140000000000000) 
14'h1ea1 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000; // D (0x00000000000000000240000000000000) 
14'h2268 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000010001000000000000000000000000000000000000000000000000000000; // D (0x00000000000000000440000000000000) 
14'h188d : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000100001000000000000000000000000000000000000000000000000000000; // D (0x00000000000000000840000000000000) 
14'h2e30 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000001000001000000000000000000000000000000000000000000000000000000; // D (0x00000000000000001040000000000000) 
14'h003d : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000010000001000000000000000000000000000000000000000000000000000000; // D (0x00000000000000002040000000000000) 
14'h1f50 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000100000001000000000000000000000000000000000000000000000000000000; // D (0x00000000000000004040000000000000) 
14'h218a : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000001000000001000000000000000000000000000000000000000000000000000000; // D (0x00000000000000008040000000000000) 
14'h1f49 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000; // D (0x00000000000000010040000000000000) 
14'h21b8 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000100000000001000000000000000000000000000000000000000000000000000000; // D (0x00000000000000020040000000000000) 
14'h1f2d : LOC =         127'b0000000000000000000000000000000000000000000000000000000000001000000000001000000000000000000000000000000000000000000000000000000; // D (0x00000000000000040040000000000000) 
14'h2170 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000010000000000001000000000000000000000000000000000000000000000000000000; // D (0x00000000000000080040000000000000) 
14'h1ebd : LOC =         127'b0000000000000000000000000000000000000000000000000000000000100000000000001000000000000000000000000000000000000000000000000000000; // D (0x00000000000000100040000000000000) 
14'h2250 : LOC =         127'b0000000000000000000000000000000000000000000000000000000001000000000000001000000000000000000000000000000000000000000000000000000; // D (0x00000000000000200040000000000000) 
14'h18fd : LOC =         127'b0000000000000000000000000000000000000000000000000000000010000000000000001000000000000000000000000000000000000000000000000000000; // D (0x00000000000000400040000000000000) 
14'h2ed0 : LOC =         127'b0000000000000000000000000000000000000000000000000000000100000000000000001000000000000000000000000000000000000000000000000000000; // D (0x00000000000000800040000000000000) 
14'h01fd : LOC =         127'b0000000000000000000000000000000000000000000000000000001000000000000000001000000000000000000000000000000000000000000000000000000; // D (0x00000000000001000040000000000000) 
14'h1cd0 : LOC =         127'b0000000000000000000000000000000000000000000000000000010000000000000000001000000000000000000000000000000000000000000000000000000; // D (0x00000000000002000040000000000000) 
14'h268a : LOC =         127'b0000000000000000000000000000000000000000000000000000100000000000000000001000000000000000000000000000000000000000000000000000000; // D (0x00000000000004000040000000000000) 
14'h1149 : LOC =         127'b0000000000000000000000000000000000000000000000000001000000000000000000001000000000000000000000000000000000000000000000000000000; // D (0x00000000000008000040000000000000) 
14'h3db8 : LOC =         127'b0000000000000000000000000000000000000000000000000010000000000000000000001000000000000000000000000000000000000000000000000000000; // D (0x00000000000010000040000000000000) 
14'h272d : LOC =         127'b0000000000000000000000000000000000000000000000000100000000000000000000001000000000000000000000000000000000000000000000000000000; // D (0x00000000000020000040000000000000) 
14'h1207 : LOC =         127'b0000000000000000000000000000000000000000000000001000000000000000000000001000000000000000000000000000000000000000000000000000000; // D (0x00000000000040000040000000000000) 
14'h3b24 : LOC =         127'b0000000000000000000000000000000000000000000000010000000000000000000000001000000000000000000000000000000000000000000000000000000; // D (0x00000000000080000040000000000000) 
14'h2a15 : LOC =         127'b0000000000000000000000000000000000000000000000100000000000000000000000001000000000000000000000000000000000000000000000000000000; // D (0x00000000000100000040000000000000) 
14'h0877 : LOC =         127'b0000000000000000000000000000000000000000000001000000000000000000000000001000000000000000000000000000000000000000000000000000000; // D (0x00000000000200000040000000000000) 
14'h0fc4 : LOC =         127'b0000000000000000000000000000000000000000000010000000000000000000000000001000000000000000000000000000000000000000000000000000000; // D (0x00000000000400000040000000000000) 
14'h00a2 : LOC =         127'b0000000000000000000000000000000000000000000100000000000000000000000000001000000000000000000000000000000000000000000000000000000; // D (0x00000000000800000040000000000000) 
14'h1e6e : LOC =         127'b0000000000000000000000000000000000000000001000000000000000000000000000001000000000000000000000000000000000000000000000000000000; // D (0x00000000001000000040000000000000) 
14'h23f6 : LOC =         127'b0000000000000000000000000000000000000000010000000000000000000000000000001000000000000000000000000000000000000000000000000000000; // D (0x00000000002000000040000000000000) 
14'h1bb1 : LOC =         127'b0000000000000000000000000000000000000000100000000000000000000000000000001000000000000000000000000000000000000000000000000000000; // D (0x00000000004000000040000000000000) 
14'h2848 : LOC =         127'b0000000000000000000000000000000000000001000000000000000000000000000000001000000000000000000000000000000000000000000000000000000; // D (0x00000000008000000040000000000000) 
14'h0ccd : LOC =         127'b0000000000000000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000000000000000000000000000; // D (0x00000000010000000040000000000000) 
14'h06b0 : LOC =         127'b0000000000000000000000000000000000000100000000000000000000000000000000001000000000000000000000000000000000000000000000000000000; // D (0x00000000020000000040000000000000) 
14'h124a : LOC =         127'b0000000000000000000000000000000000001000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000; // D (0x00000000040000000040000000000000) 
14'h3bbe : LOC =         127'b0000000000000000000000000000000000010000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000; // D (0x00000000080000000040000000000000) 
14'h2b21 : LOC =         127'b0000000000000000000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000; // D (0x00000000100000000040000000000000) 
14'h0a1f : LOC =         127'b0000000000000000000000000000000001000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000; // D (0x00000000200000000040000000000000) 
14'h0b14 : LOC =         127'b0000000000000000000000000000000010000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000; // D (0x00000000400000000040000000000000) 
14'h0902 : LOC =         127'b0000000000000000000000000000000100000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000; // D (0x00000000800000000040000000000000) 
14'h0d2e : LOC =         127'b0000000000000000000000000000001000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000; // D (0x00000001000000000040000000000000) 
14'h0576 : LOC =         127'b0000000000000000000000000000010000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000; // D (0x00000002000000000040000000000000) 
14'h15c6 : LOC =         127'b0000000000000000000000000000100000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000; // D (0x00000004000000000040000000000000) 
14'h34a6 : LOC =         127'b0000000000000000000000000001000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000; // D (0x00000008000000000040000000000000) 
14'h3511 : LOC =         127'b0000000000000000000000000010000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000; // D (0x00000010000000000040000000000000) 
14'h367f : LOC =         127'b0000000000000000000000000100000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000; // D (0x00000020000000000040000000000000) 
14'h30a3 : LOC =         127'b0000000000000000000000001000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000; // D (0x00000040000000000040000000000000) 
14'h3d1b : LOC =         127'b0000000000000000000000010000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000; // D (0x00000080000000000040000000000000) 
14'h266b : LOC =         127'b0000000000000000000000100000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000; // D (0x00000100000000000040000000000000) 
14'h108b : LOC =         127'b0000000000000000000001000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000; // D (0x00000200000000000040000000000000) 
14'h3e3c : LOC =         127'b0000000000000000000010000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000; // D (0x00000400000000000040000000000000) 
14'h2025 : LOC =         127'b0000000000000000000100000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000; // D (0x00000800000000000040000000000000) 
14'h1c17 : LOC =         127'b0000000000000000001000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000; // D (0x00001000000000000040000000000000) 
14'h2704 : LOC =         127'b0000000000000000010000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000; // D (0x00002000000000000040000000000000) 
14'h1255 : LOC =         127'b0000000000000000100000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000; // D (0x00004000000000000040000000000000) 
14'h3b80 : LOC =         127'b0000000000000001000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000; // D (0x00008000000000000040000000000000) 
14'h2b5d : LOC =         127'b0000000000000010000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000; // D (0x00010000000000000040000000000000) 
14'h0ae7 : LOC =         127'b0000000000000100000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000; // D (0x00020000000000000040000000000000) 
14'h0ae4 : LOC =         127'b0000000000001000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000; // D (0x00040000000000000040000000000000) 
14'h0ae2 : LOC =         127'b0000000000010000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000; // D (0x00080000000000000040000000000000) 
14'h0aee : LOC =         127'b0000000000100000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000; // D (0x00100000000000000040000000000000) 
14'h0af6 : LOC =         127'b0000000001000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000; // D (0x00200000000000000040000000000000) 
14'h0ac6 : LOC =         127'b0000000010000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000; // D (0x00400000000000000040000000000000) 
14'h0aa6 : LOC =         127'b0000000100000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000; // D (0x00800000000000000040000000000000) 
14'h0a66 : LOC =         127'b0000001000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000; // D (0x01000000000000000040000000000000) 
14'h0be6 : LOC =         127'b0000010000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000; // D (0x02000000000000000040000000000000) 
14'h08e6 : LOC =         127'b0000100000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000; // D (0x04000000000000000040000000000000) 
14'h0ee6 : LOC =         127'b0001000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000; // D (0x08000000000000000040000000000000) 
14'h02e6 : LOC =         127'b0010000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000; // D (0x10000000000000000040000000000000) 
14'h1ae6 : LOC =         127'b0100000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000; // D (0x20000000000000000040000000000000) 
14'h2ae6 : LOC =         127'b1000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000; // D (0x40000000000000000040000000000000) 
14'h15cc : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000; // S (0x00000000000000000080000000000000) 
14'h3e54 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000000000000000000000000000000000000; // D (0x00000000000000000180000000000000) 
14'h018b : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000001010000000000000000000000000000000000000000000000000000000; // D (0x00000000000000000280000000000000) 
14'h3d42 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000; // D (0x00000000000000000480000000000000) 
14'h07a7 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000100010000000000000000000000000000000000000000000000000000000; // D (0x00000000000000000880000000000000) 
14'h311a : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000001000010000000000000000000000000000000000000000000000000000000; // D (0x00000000000000001080000000000000) 
14'h1f17 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000010000010000000000000000000000000000000000000000000000000000000; // D (0x00000000000000002080000000000000) 
14'h007a : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000100000010000000000000000000000000000000000000000000000000000000; // D (0x00000000000000004080000000000000) 
14'h3ea0 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000001000000010000000000000000000000000000000000000000000000000000000; // D (0x00000000000000008080000000000000) 
14'h0063 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000010000000010000000000000000000000000000000000000000000000000000000; // D (0x00000000000000010080000000000000) 
14'h3e92 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000100000000010000000000000000000000000000000000000000000000000000000; // D (0x00000000000000020080000000000000) 
14'h0007 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000001000000000010000000000000000000000000000000000000000000000000000000; // D (0x00000000000000040080000000000000) 
14'h3e5a : LOC =         127'b0000000000000000000000000000000000000000000000000000000000010000000000010000000000000000000000000000000000000000000000000000000; // D (0x00000000000000080080000000000000) 
14'h0197 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000100000000000010000000000000000000000000000000000000000000000000000000; // D (0x00000000000000100080000000000000) 
14'h3d7a : LOC =         127'b0000000000000000000000000000000000000000000000000000000001000000000000010000000000000000000000000000000000000000000000000000000; // D (0x00000000000000200080000000000000) 
14'h07d7 : LOC =         127'b0000000000000000000000000000000000000000000000000000000010000000000000010000000000000000000000000000000000000000000000000000000; // D (0x00000000000000400080000000000000) 
14'h31fa : LOC =         127'b0000000000000000000000000000000000000000000000000000000100000000000000010000000000000000000000000000000000000000000000000000000; // D (0x00000000000000800080000000000000) 
14'h1ed7 : LOC =         127'b0000000000000000000000000000000000000000000000000000001000000000000000010000000000000000000000000000000000000000000000000000000; // D (0x00000000000001000080000000000000) 
14'h03fa : LOC =         127'b0000000000000000000000000000000000000000000000000000010000000000000000010000000000000000000000000000000000000000000000000000000; // D (0x00000000000002000080000000000000) 
14'h39a0 : LOC =         127'b0000000000000000000000000000000000000000000000000000100000000000000000010000000000000000000000000000000000000000000000000000000; // D (0x00000000000004000080000000000000) 
14'h0e63 : LOC =         127'b0000000000000000000000000000000000000000000000000001000000000000000000010000000000000000000000000000000000000000000000000000000; // D (0x00000000000008000080000000000000) 
14'h2292 : LOC =         127'b0000000000000000000000000000000000000000000000000010000000000000000000010000000000000000000000000000000000000000000000000000000; // D (0x00000000000010000080000000000000) 
14'h3807 : LOC =         127'b0000000000000000000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000000000000000000000000; // D (0x00000000000020000080000000000000) 
14'h0d2d : LOC =         127'b0000000000000000000000000000000000000000000000001000000000000000000000010000000000000000000000000000000000000000000000000000000; // D (0x00000000000040000080000000000000) 
14'h240e : LOC =         127'b0000000000000000000000000000000000000000000000010000000000000000000000010000000000000000000000000000000000000000000000000000000; // D (0x00000000000080000080000000000000) 
14'h353f : LOC =         127'b0000000000000000000000000000000000000000000000100000000000000000000000010000000000000000000000000000000000000000000000000000000; // D (0x00000000000100000080000000000000) 
14'h175d : LOC =         127'b0000000000000000000000000000000000000000000001000000000000000000000000010000000000000000000000000000000000000000000000000000000; // D (0x00000000000200000080000000000000) 
14'h10ee : LOC =         127'b0000000000000000000000000000000000000000000010000000000000000000000000010000000000000000000000000000000000000000000000000000000; // D (0x00000000000400000080000000000000) 
14'h1f88 : LOC =         127'b0000000000000000000000000000000000000000000100000000000000000000000000010000000000000000000000000000000000000000000000000000000; // D (0x00000000000800000080000000000000) 
14'h0144 : LOC =         127'b0000000000000000000000000000000000000000001000000000000000000000000000010000000000000000000000000000000000000000000000000000000; // D (0x00000000001000000080000000000000) 
14'h3cdc : LOC =         127'b0000000000000000000000000000000000000000010000000000000000000000000000010000000000000000000000000000000000000000000000000000000; // D (0x00000000002000000080000000000000) 
14'h049b : LOC =         127'b0000000000000000000000000000000000000000100000000000000000000000000000010000000000000000000000000000000000000000000000000000000; // D (0x00000000004000000080000000000000) 
14'h3762 : LOC =         127'b0000000000000000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000000000000000000000000000; // D (0x00000000008000000080000000000000) 
14'h13e7 : LOC =         127'b0000000000000000000000000000000000000010000000000000000000000000000000010000000000000000000000000000000000000000000000000000000; // D (0x00000000010000000080000000000000) 
14'h199a : LOC =         127'b0000000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000000000000000000000000; // D (0x00000000020000000080000000000000) 
14'h0d60 : LOC =         127'b0000000000000000000000000000000000001000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000; // D (0x00000000040000000080000000000000) 
14'h2494 : LOC =         127'b0000000000000000000000000000000000010000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000; // D (0x00000000080000000080000000000000) 
14'h340b : LOC =         127'b0000000000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000; // D (0x00000000100000000080000000000000) 
14'h1535 : LOC =         127'b0000000000000000000000000000000001000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000; // D (0x00000000200000000080000000000000) 
14'h143e : LOC =         127'b0000000000000000000000000000000010000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000; // D (0x00000000400000000080000000000000) 
14'h1628 : LOC =         127'b0000000000000000000000000000000100000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000; // D (0x00000000800000000080000000000000) 
14'h1204 : LOC =         127'b0000000000000000000000000000001000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000; // D (0x00000001000000000080000000000000) 
14'h1a5c : LOC =         127'b0000000000000000000000000000010000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000; // D (0x00000002000000000080000000000000) 
14'h0aec : LOC =         127'b0000000000000000000000000000100000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000; // D (0x00000004000000000080000000000000) 
14'h2b8c : LOC =         127'b0000000000000000000000000001000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000; // D (0x00000008000000000080000000000000) 
14'h2a3b : LOC =         127'b0000000000000000000000000010000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000; // D (0x00000010000000000080000000000000) 
14'h2955 : LOC =         127'b0000000000000000000000000100000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000; // D (0x00000020000000000080000000000000) 
14'h2f89 : LOC =         127'b0000000000000000000000001000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000; // D (0x00000040000000000080000000000000) 
14'h2231 : LOC =         127'b0000000000000000000000010000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000; // D (0x00000080000000000080000000000000) 
14'h3941 : LOC =         127'b0000000000000000000000100000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000; // D (0x00000100000000000080000000000000) 
14'h0fa1 : LOC =         127'b0000000000000000000001000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000; // D (0x00000200000000000080000000000000) 
14'h2116 : LOC =         127'b0000000000000000000010000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000; // D (0x00000400000000000080000000000000) 
14'h3f0f : LOC =         127'b0000000000000000000100000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000; // D (0x00000800000000000080000000000000) 
14'h033d : LOC =         127'b0000000000000000001000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000; // D (0x00001000000000000080000000000000) 
14'h382e : LOC =         127'b0000000000000000010000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000; // D (0x00002000000000000080000000000000) 
14'h0d7f : LOC =         127'b0000000000000000100000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000; // D (0x00004000000000000080000000000000) 
14'h24aa : LOC =         127'b0000000000000001000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000; // D (0x00008000000000000080000000000000) 
14'h3477 : LOC =         127'b0000000000000010000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000; // D (0x00010000000000000080000000000000) 
14'h15cd : LOC =         127'b0000000000000100000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000; // D (0x00020000000000000080000000000000) 
14'h15ce : LOC =         127'b0000000000001000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000; // D (0x00040000000000000080000000000000) 
14'h15c8 : LOC =         127'b0000000000010000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000; // D (0x00080000000000000080000000000000) 
14'h15c4 : LOC =         127'b0000000000100000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000; // D (0x00100000000000000080000000000000) 
14'h15dc : LOC =         127'b0000000001000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000; // D (0x00200000000000000080000000000000) 
14'h15ec : LOC =         127'b0000000010000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000; // D (0x00400000000000000080000000000000) 
14'h158c : LOC =         127'b0000000100000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000; // D (0x00800000000000000080000000000000) 
14'h154c : LOC =         127'b0000001000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000; // D (0x01000000000000000080000000000000) 
14'h14cc : LOC =         127'b0000010000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000; // D (0x02000000000000000080000000000000) 
14'h17cc : LOC =         127'b0000100000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000; // D (0x04000000000000000080000000000000) 
14'h11cc : LOC =         127'b0001000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000; // D (0x08000000000000000080000000000000) 
14'h1dcc : LOC =         127'b0010000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000; // D (0x10000000000000000080000000000000) 
14'h05cc : LOC =         127'b0100000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000; // D (0x20000000000000000080000000000000) 
14'h35cc : LOC =         127'b1000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000; // D (0x40000000000000000080000000000000) 
14'h2b98 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000; // S (0x00000000000000000100000000000000) 
14'h3fdf : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000; // D (0x00000000000000000300000000000000) 
14'h0316 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000000000000000000000000000000000; // D (0x00000000000000000500000000000000) 
14'h39f3 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000; // D (0x00000000000000000900000000000000) 
14'h0f4e : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000001000100000000000000000000000000000000000000000000000000000000; // D (0x00000000000000001100000000000000) 
14'h2143 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000010000100000000000000000000000000000000000000000000000000000000; // D (0x00000000000000002100000000000000) 
14'h3e2e : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000100000100000000000000000000000000000000000000000000000000000000; // D (0x00000000000000004100000000000000) 
14'h00f4 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000001000000100000000000000000000000000000000000000000000000000000000; // D (0x00000000000000008100000000000000) 
14'h3e37 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000010000000100000000000000000000000000000000000000000000000000000000; // D (0x00000000000000010100000000000000) 
14'h00c6 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000100000000100000000000000000000000000000000000000000000000000000000; // D (0x00000000000000020100000000000000) 
14'h3e53 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000001000000000100000000000000000000000000000000000000000000000000000000; // D (0x00000000000000040100000000000000) 
14'h000e : LOC =         127'b0000000000000000000000000000000000000000000000000000000000010000000000100000000000000000000000000000000000000000000000000000000; // D (0x00000000000000080100000000000000) 
14'h3fc3 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000100000000000100000000000000000000000000000000000000000000000000000000; // D (0x00000000000000100100000000000000) 
14'h032e : LOC =         127'b0000000000000000000000000000000000000000000000000000000001000000000000100000000000000000000000000000000000000000000000000000000; // D (0x00000000000000200100000000000000) 
14'h3983 : LOC =         127'b0000000000000000000000000000000000000000000000000000000010000000000000100000000000000000000000000000000000000000000000000000000; // D (0x00000000000000400100000000000000) 
14'h0fae : LOC =         127'b0000000000000000000000000000000000000000000000000000000100000000000000100000000000000000000000000000000000000000000000000000000; // D (0x00000000000000800100000000000000) 
14'h2083 : LOC =         127'b0000000000000000000000000000000000000000000000000000001000000000000000100000000000000000000000000000000000000000000000000000000; // D (0x00000000000001000100000000000000) 
14'h3dae : LOC =         127'b0000000000000000000000000000000000000000000000000000010000000000000000100000000000000000000000000000000000000000000000000000000; // D (0x00000000000002000100000000000000) 
14'h07f4 : LOC =         127'b0000000000000000000000000000000000000000000000000000100000000000000000100000000000000000000000000000000000000000000000000000000; // D (0x00000000000004000100000000000000) 
14'h3037 : LOC =         127'b0000000000000000000000000000000000000000000000000001000000000000000000100000000000000000000000000000000000000000000000000000000; // D (0x00000000000008000100000000000000) 
14'h1cc6 : LOC =         127'b0000000000000000000000000000000000000000000000000010000000000000000000100000000000000000000000000000000000000000000000000000000; // D (0x00000000000010000100000000000000) 
14'h0653 : LOC =         127'b0000000000000000000000000000000000000000000000000100000000000000000000100000000000000000000000000000000000000000000000000000000; // D (0x00000000000020000100000000000000) 
14'h3379 : LOC =         127'b0000000000000000000000000000000000000000000000001000000000000000000000100000000000000000000000000000000000000000000000000000000; // D (0x00000000000040000100000000000000) 
14'h1a5a : LOC =         127'b0000000000000000000000000000000000000000000000010000000000000000000000100000000000000000000000000000000000000000000000000000000; // D (0x00000000000080000100000000000000) 
14'h0b6b : LOC =         127'b0000000000000000000000000000000000000000000000100000000000000000000000100000000000000000000000000000000000000000000000000000000; // D (0x00000000000100000100000000000000) 
14'h2909 : LOC =         127'b0000000000000000000000000000000000000000000001000000000000000000000000100000000000000000000000000000000000000000000000000000000; // D (0x00000000000200000100000000000000) 
14'h2eba : LOC =         127'b0000000000000000000000000000000000000000000010000000000000000000000000100000000000000000000000000000000000000000000000000000000; // D (0x00000000000400000100000000000000) 
14'h21dc : LOC =         127'b0000000000000000000000000000000000000000000100000000000000000000000000100000000000000000000000000000000000000000000000000000000; // D (0x00000000000800000100000000000000) 
14'h3f10 : LOC =         127'b0000000000000000000000000000000000000000001000000000000000000000000000100000000000000000000000000000000000000000000000000000000; // D (0x00000000001000000100000000000000) 
14'h0288 : LOC =         127'b0000000000000000000000000000000000000000010000000000000000000000000000100000000000000000000000000000000000000000000000000000000; // D (0x00000000002000000100000000000000) 
14'h3acf : LOC =         127'b0000000000000000000000000000000000000000100000000000000000000000000000100000000000000000000000000000000000000000000000000000000; // D (0x00000000004000000100000000000000) 
14'h0936 : LOC =         127'b0000000000000000000000000000000000000001000000000000000000000000000000100000000000000000000000000000000000000000000000000000000; // D (0x00000000008000000100000000000000) 
14'h2db3 : LOC =         127'b0000000000000000000000000000000000000010000000000000000000000000000000100000000000000000000000000000000000000000000000000000000; // D (0x00000000010000000100000000000000) 
14'h27ce : LOC =         127'b0000000000000000000000000000000000000100000000000000000000000000000000100000000000000000000000000000000000000000000000000000000; // D (0x00000000020000000100000000000000) 
14'h3334 : LOC =         127'b0000000000000000000000000000000000001000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000; // D (0x00000000040000000100000000000000) 
14'h1ac0 : LOC =         127'b0000000000000000000000000000000000010000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000; // D (0x00000000080000000100000000000000) 
14'h0a5f : LOC =         127'b0000000000000000000000000000000000100000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000; // D (0x00000000100000000100000000000000) 
14'h2b61 : LOC =         127'b0000000000000000000000000000000001000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000; // D (0x00000000200000000100000000000000) 
14'h2a6a : LOC =         127'b0000000000000000000000000000000010000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000; // D (0x00000000400000000100000000000000) 
14'h287c : LOC =         127'b0000000000000000000000000000000100000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000; // D (0x00000000800000000100000000000000) 
14'h2c50 : LOC =         127'b0000000000000000000000000000001000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000; // D (0x00000001000000000100000000000000) 
14'h2408 : LOC =         127'b0000000000000000000000000000010000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000; // D (0x00000002000000000100000000000000) 
14'h34b8 : LOC =         127'b0000000000000000000000000000100000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000; // D (0x00000004000000000100000000000000) 
14'h15d8 : LOC =         127'b0000000000000000000000000001000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000; // D (0x00000008000000000100000000000000) 
14'h146f : LOC =         127'b0000000000000000000000000010000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000; // D (0x00000010000000000100000000000000) 
14'h1701 : LOC =         127'b0000000000000000000000000100000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000; // D (0x00000020000000000100000000000000) 
14'h11dd : LOC =         127'b0000000000000000000000001000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000; // D (0x00000040000000000100000000000000) 
14'h1c65 : LOC =         127'b0000000000000000000000010000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000; // D (0x00000080000000000100000000000000) 
14'h0715 : LOC =         127'b0000000000000000000000100000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000; // D (0x00000100000000000100000000000000) 
14'h31f5 : LOC =         127'b0000000000000000000001000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000; // D (0x00000200000000000100000000000000) 
14'h1f42 : LOC =         127'b0000000000000000000010000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000; // D (0x00000400000000000100000000000000) 
14'h015b : LOC =         127'b0000000000000000000100000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000; // D (0x00000800000000000100000000000000) 
14'h3d69 : LOC =         127'b0000000000000000001000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000; // D (0x00001000000000000100000000000000) 
14'h067a : LOC =         127'b0000000000000000010000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000; // D (0x00002000000000000100000000000000) 
14'h332b : LOC =         127'b0000000000000000100000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000; // D (0x00004000000000000100000000000000) 
14'h1afe : LOC =         127'b0000000000000001000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000; // D (0x00008000000000000100000000000000) 
14'h0a23 : LOC =         127'b0000000000000010000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000; // D (0x00010000000000000100000000000000) 
14'h2b99 : LOC =         127'b0000000000000100000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000; // D (0x00020000000000000100000000000000) 
14'h2b9a : LOC =         127'b0000000000001000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000; // D (0x00040000000000000100000000000000) 
14'h2b9c : LOC =         127'b0000000000010000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000; // D (0x00080000000000000100000000000000) 
14'h2b90 : LOC =         127'b0000000000100000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000; // D (0x00100000000000000100000000000000) 
14'h2b88 : LOC =         127'b0000000001000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000; // D (0x00200000000000000100000000000000) 
14'h2bb8 : LOC =         127'b0000000010000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000; // D (0x00400000000000000100000000000000) 
14'h2bd8 : LOC =         127'b0000000100000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000; // D (0x00800000000000000100000000000000) 
14'h2b18 : LOC =         127'b0000001000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000; // D (0x01000000000000000100000000000000) 
14'h2a98 : LOC =         127'b0000010000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000; // D (0x02000000000000000100000000000000) 
14'h2998 : LOC =         127'b0000100000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000; // D (0x04000000000000000100000000000000) 
14'h2f98 : LOC =         127'b0001000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000; // D (0x08000000000000000100000000000000) 
14'h2398 : LOC =         127'b0010000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000; // D (0x10000000000000000100000000000000) 
14'h3b98 : LOC =         127'b0100000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000; // D (0x20000000000000000100000000000000) 
14'h0b98 : LOC =         127'b1000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000; // D (0x40000000000000000100000000000000) 
14'h1447 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000; // S (0x00000000000000000200000000000000) 
14'h3cc9 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000000000000000000000000000000000000; // D (0x00000000000000000600000000000000) 
14'h062c : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000101000000000000000000000000000000000000000000000000000000000; // D (0x00000000000000000a00000000000000) 
14'h3091 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000; // D (0x00000000000000001200000000000000) 
14'h1e9c : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000010001000000000000000000000000000000000000000000000000000000000; // D (0x00000000000000002200000000000000) 
14'h01f1 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000100001000000000000000000000000000000000000000000000000000000000; // D (0x00000000000000004200000000000000) 
14'h3f2b : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000001000001000000000000000000000000000000000000000000000000000000000; // D (0x00000000000000008200000000000000) 
14'h01e8 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000010000001000000000000000000000000000000000000000000000000000000000; // D (0x00000000000000010200000000000000) 
14'h3f19 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000100000001000000000000000000000000000000000000000000000000000000000; // D (0x00000000000000020200000000000000) 
14'h018c : LOC =         127'b0000000000000000000000000000000000000000000000000000000000001000000001000000000000000000000000000000000000000000000000000000000; // D (0x00000000000000040200000000000000) 
14'h3fd1 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000000; // D (0x00000000000000080200000000000000) 
14'h001c : LOC =         127'b0000000000000000000000000000000000000000000000000000000000100000000001000000000000000000000000000000000000000000000000000000000; // D (0x00000000000000100200000000000000) 
14'h3cf1 : LOC =         127'b0000000000000000000000000000000000000000000000000000000001000000000001000000000000000000000000000000000000000000000000000000000; // D (0x00000000000000200200000000000000) 
14'h065c : LOC =         127'b0000000000000000000000000000000000000000000000000000000010000000000001000000000000000000000000000000000000000000000000000000000; // D (0x00000000000000400200000000000000) 
14'h3071 : LOC =         127'b0000000000000000000000000000000000000000000000000000000100000000000001000000000000000000000000000000000000000000000000000000000; // D (0x00000000000000800200000000000000) 
14'h1f5c : LOC =         127'b0000000000000000000000000000000000000000000000000000001000000000000001000000000000000000000000000000000000000000000000000000000; // D (0x00000000000001000200000000000000) 
14'h0271 : LOC =         127'b0000000000000000000000000000000000000000000000000000010000000000000001000000000000000000000000000000000000000000000000000000000; // D (0x00000000000002000200000000000000) 
14'h382b : LOC =         127'b0000000000000000000000000000000000000000000000000000100000000000000001000000000000000000000000000000000000000000000000000000000; // D (0x00000000000004000200000000000000) 
14'h0fe8 : LOC =         127'b0000000000000000000000000000000000000000000000000001000000000000000001000000000000000000000000000000000000000000000000000000000; // D (0x00000000000008000200000000000000) 
14'h2319 : LOC =         127'b0000000000000000000000000000000000000000000000000010000000000000000001000000000000000000000000000000000000000000000000000000000; // D (0x00000000000010000200000000000000) 
14'h398c : LOC =         127'b0000000000000000000000000000000000000000000000000100000000000000000001000000000000000000000000000000000000000000000000000000000; // D (0x00000000000020000200000000000000) 
14'h0ca6 : LOC =         127'b0000000000000000000000000000000000000000000000001000000000000000000001000000000000000000000000000000000000000000000000000000000; // D (0x00000000000040000200000000000000) 
14'h2585 : LOC =         127'b0000000000000000000000000000000000000000000000010000000000000000000001000000000000000000000000000000000000000000000000000000000; // D (0x00000000000080000200000000000000) 
14'h34b4 : LOC =         127'b0000000000000000000000000000000000000000000000100000000000000000000001000000000000000000000000000000000000000000000000000000000; // D (0x00000000000100000200000000000000) 
14'h16d6 : LOC =         127'b0000000000000000000000000000000000000000000001000000000000000000000001000000000000000000000000000000000000000000000000000000000; // D (0x00000000000200000200000000000000) 
14'h1165 : LOC =         127'b0000000000000000000000000000000000000000000010000000000000000000000001000000000000000000000000000000000000000000000000000000000; // D (0x00000000000400000200000000000000) 
14'h1e03 : LOC =         127'b0000000000000000000000000000000000000000000100000000000000000000000001000000000000000000000000000000000000000000000000000000000; // D (0x00000000000800000200000000000000) 
14'h00cf : LOC =         127'b0000000000000000000000000000000000000000001000000000000000000000000001000000000000000000000000000000000000000000000000000000000; // D (0x00000000001000000200000000000000) 
14'h3d57 : LOC =         127'b0000000000000000000000000000000000000000010000000000000000000000000001000000000000000000000000000000000000000000000000000000000; // D (0x00000000002000000200000000000000) 
14'h0510 : LOC =         127'b0000000000000000000000000000000000000000100000000000000000000000000001000000000000000000000000000000000000000000000000000000000; // D (0x00000000004000000200000000000000) 
14'h36e9 : LOC =         127'b0000000000000000000000000000000000000001000000000000000000000000000001000000000000000000000000000000000000000000000000000000000; // D (0x00000000008000000200000000000000) 
14'h126c : LOC =         127'b0000000000000000000000000000000000000010000000000000000000000000000001000000000000000000000000000000000000000000000000000000000; // D (0x00000000010000000200000000000000) 
14'h1811 : LOC =         127'b0000000000000000000000000000000000000100000000000000000000000000000001000000000000000000000000000000000000000000000000000000000; // D (0x00000000020000000200000000000000) 
14'h0ceb : LOC =         127'b0000000000000000000000000000000000001000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000; // D (0x00000000040000000200000000000000) 
14'h251f : LOC =         127'b0000000000000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000; // D (0x00000000080000000200000000000000) 
14'h3580 : LOC =         127'b0000000000000000000000000000000000100000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000; // D (0x00000000100000000200000000000000) 
14'h14be : LOC =         127'b0000000000000000000000000000000001000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000; // D (0x00000000200000000200000000000000) 
14'h15b5 : LOC =         127'b0000000000000000000000000000000010000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000; // D (0x00000000400000000200000000000000) 
14'h17a3 : LOC =         127'b0000000000000000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000; // D (0x00000000800000000200000000000000) 
14'h138f : LOC =         127'b0000000000000000000000000000001000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000; // D (0x00000001000000000200000000000000) 
14'h1bd7 : LOC =         127'b0000000000000000000000000000010000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000; // D (0x00000002000000000200000000000000) 
14'h0b67 : LOC =         127'b0000000000000000000000000000100000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000; // D (0x00000004000000000200000000000000) 
14'h2a07 : LOC =         127'b0000000000000000000000000001000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000; // D (0x00000008000000000200000000000000) 
14'h2bb0 : LOC =         127'b0000000000000000000000000010000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000; // D (0x00000010000000000200000000000000) 
14'h28de : LOC =         127'b0000000000000000000000000100000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000; // D (0x00000020000000000200000000000000) 
14'h2e02 : LOC =         127'b0000000000000000000000001000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000; // D (0x00000040000000000200000000000000) 
14'h23ba : LOC =         127'b0000000000000000000000010000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000; // D (0x00000080000000000200000000000000) 
14'h38ca : LOC =         127'b0000000000000000000000100000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000; // D (0x00000100000000000200000000000000) 
14'h0e2a : LOC =         127'b0000000000000000000001000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000; // D (0x00000200000000000200000000000000) 
14'h209d : LOC =         127'b0000000000000000000010000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000; // D (0x00000400000000000200000000000000) 
14'h3e84 : LOC =         127'b0000000000000000000100000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000; // D (0x00000800000000000200000000000000) 
14'h02b6 : LOC =         127'b0000000000000000001000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000; // D (0x00001000000000000200000000000000) 
14'h39a5 : LOC =         127'b0000000000000000010000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000; // D (0x00002000000000000200000000000000) 
14'h0cf4 : LOC =         127'b0000000000000000100000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000; // D (0x00004000000000000200000000000000) 
14'h2521 : LOC =         127'b0000000000000001000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000; // D (0x00008000000000000200000000000000) 
14'h35fc : LOC =         127'b0000000000000010000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000; // D (0x00010000000000000200000000000000) 
14'h1446 : LOC =         127'b0000000000000100000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000; // D (0x00020000000000000200000000000000) 
14'h1445 : LOC =         127'b0000000000001000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000; // D (0x00040000000000000200000000000000) 
14'h1443 : LOC =         127'b0000000000010000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000; // D (0x00080000000000000200000000000000) 
14'h144f : LOC =         127'b0000000000100000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000; // D (0x00100000000000000200000000000000) 
14'h1457 : LOC =         127'b0000000001000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000; // D (0x00200000000000000200000000000000) 
14'h1467 : LOC =         127'b0000000010000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000; // D (0x00400000000000000200000000000000) 
14'h1407 : LOC =         127'b0000000100000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000; // D (0x00800000000000000200000000000000) 
14'h14c7 : LOC =         127'b0000001000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000; // D (0x01000000000000000200000000000000) 
14'h1547 : LOC =         127'b0000010000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000; // D (0x02000000000000000200000000000000) 
14'h1647 : LOC =         127'b0000100000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000; // D (0x04000000000000000200000000000000) 
14'h1047 : LOC =         127'b0001000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000; // D (0x08000000000000000200000000000000) 
14'h1c47 : LOC =         127'b0010000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000; // D (0x10000000000000000200000000000000) 
14'h0447 : LOC =         127'b0100000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000; // D (0x20000000000000000200000000000000) 
14'h3447 : LOC =         127'b1000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000; // D (0x40000000000000000200000000000000) 
14'h288e : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000; // S (0x00000000000000000400000000000000) 
14'h3ae5 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000; // D (0x00000000000000000c00000000000000) 
14'h0c58 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000001010000000000000000000000000000000000000000000000000000000000; // D (0x00000000000000001400000000000000) 
14'h2255 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000; // D (0x00000000000000002400000000000000) 
14'h3d38 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000100010000000000000000000000000000000000000000000000000000000000; // D (0x00000000000000004400000000000000) 
14'h03e2 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000001000010000000000000000000000000000000000000000000000000000000000; // D (0x00000000000000008400000000000000) 
14'h3d21 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000010000010000000000000000000000000000000000000000000000000000000000; // D (0x00000000000000010400000000000000) 
14'h03d0 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000100000010000000000000000000000000000000000000000000000000000000000; // D (0x00000000000000020400000000000000) 
14'h3d45 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000001000000010000000000000000000000000000000000000000000000000000000000; // D (0x00000000000000040400000000000000) 
14'h0318 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000010000000010000000000000000000000000000000000000000000000000000000000; // D (0x00000000000000080400000000000000) 
14'h3cd5 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000100000000010000000000000000000000000000000000000000000000000000000000; // D (0x00000000000000100400000000000000) 
14'h0038 : LOC =         127'b0000000000000000000000000000000000000000000000000000000001000000000010000000000000000000000000000000000000000000000000000000000; // D (0x00000000000000200400000000000000) 
14'h3a95 : LOC =         127'b0000000000000000000000000000000000000000000000000000000010000000000010000000000000000000000000000000000000000000000000000000000; // D (0x00000000000000400400000000000000) 
14'h0cb8 : LOC =         127'b0000000000000000000000000000000000000000000000000000000100000000000010000000000000000000000000000000000000000000000000000000000; // D (0x00000000000000800400000000000000) 
14'h2395 : LOC =         127'b0000000000000000000000000000000000000000000000000000001000000000000010000000000000000000000000000000000000000000000000000000000; // D (0x00000000000001000400000000000000) 
14'h3eb8 : LOC =         127'b0000000000000000000000000000000000000000000000000000010000000000000010000000000000000000000000000000000000000000000000000000000; // D (0x00000000000002000400000000000000) 
14'h04e2 : LOC =         127'b0000000000000000000000000000000000000000000000000000100000000000000010000000000000000000000000000000000000000000000000000000000; // D (0x00000000000004000400000000000000) 
14'h3321 : LOC =         127'b0000000000000000000000000000000000000000000000000001000000000000000010000000000000000000000000000000000000000000000000000000000; // D (0x00000000000008000400000000000000) 
14'h1fd0 : LOC =         127'b0000000000000000000000000000000000000000000000000010000000000000000010000000000000000000000000000000000000000000000000000000000; // D (0x00000000000010000400000000000000) 
14'h0545 : LOC =         127'b0000000000000000000000000000000000000000000000000100000000000000000010000000000000000000000000000000000000000000000000000000000; // D (0x00000000000020000400000000000000) 
14'h306f : LOC =         127'b0000000000000000000000000000000000000000000000001000000000000000000010000000000000000000000000000000000000000000000000000000000; // D (0x00000000000040000400000000000000) 
14'h194c : LOC =         127'b0000000000000000000000000000000000000000000000010000000000000000000010000000000000000000000000000000000000000000000000000000000; // D (0x00000000000080000400000000000000) 
14'h087d : LOC =         127'b0000000000000000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000000000000000000000000000; // D (0x00000000000100000400000000000000) 
14'h2a1f : LOC =         127'b0000000000000000000000000000000000000000000001000000000000000000000010000000000000000000000000000000000000000000000000000000000; // D (0x00000000000200000400000000000000) 
14'h2dac : LOC =         127'b0000000000000000000000000000000000000000000010000000000000000000000010000000000000000000000000000000000000000000000000000000000; // D (0x00000000000400000400000000000000) 
14'h22ca : LOC =         127'b0000000000000000000000000000000000000000000100000000000000000000000010000000000000000000000000000000000000000000000000000000000; // D (0x00000000000800000400000000000000) 
14'h3c06 : LOC =         127'b0000000000000000000000000000000000000000001000000000000000000000000010000000000000000000000000000000000000000000000000000000000; // D (0x00000000001000000400000000000000) 
14'h019e : LOC =         127'b0000000000000000000000000000000000000000010000000000000000000000000010000000000000000000000000000000000000000000000000000000000; // D (0x00000000002000000400000000000000) 
14'h39d9 : LOC =         127'b0000000000000000000000000000000000000000100000000000000000000000000010000000000000000000000000000000000000000000000000000000000; // D (0x00000000004000000400000000000000) 
14'h0a20 : LOC =         127'b0000000000000000000000000000000000000001000000000000000000000000000010000000000000000000000000000000000000000000000000000000000; // D (0x00000000008000000400000000000000) 
14'h2ea5 : LOC =         127'b0000000000000000000000000000000000000010000000000000000000000000000010000000000000000000000000000000000000000000000000000000000; // D (0x00000000010000000400000000000000) 
14'h24d8 : LOC =         127'b0000000000000000000000000000000000000100000000000000000000000000000010000000000000000000000000000000000000000000000000000000000; // D (0x00000000020000000400000000000000) 
14'h3022 : LOC =         127'b0000000000000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000; // D (0x00000000040000000400000000000000) 
14'h19d6 : LOC =         127'b0000000000000000000000000000000000010000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000; // D (0x00000000080000000400000000000000) 
14'h0949 : LOC =         127'b0000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000; // D (0x00000000100000000400000000000000) 
14'h2877 : LOC =         127'b0000000000000000000000000000000001000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000; // D (0x00000000200000000400000000000000) 
14'h297c : LOC =         127'b0000000000000000000000000000000010000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000; // D (0x00000000400000000400000000000000) 
14'h2b6a : LOC =         127'b0000000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000; // D (0x00000000800000000400000000000000) 
14'h2f46 : LOC =         127'b0000000000000000000000000000001000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000; // D (0x00000001000000000400000000000000) 
14'h271e : LOC =         127'b0000000000000000000000000000010000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000; // D (0x00000002000000000400000000000000) 
14'h37ae : LOC =         127'b0000000000000000000000000000100000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000; // D (0x00000004000000000400000000000000) 
14'h16ce : LOC =         127'b0000000000000000000000000001000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000; // D (0x00000008000000000400000000000000) 
14'h1779 : LOC =         127'b0000000000000000000000000010000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000; // D (0x00000010000000000400000000000000) 
14'h1417 : LOC =         127'b0000000000000000000000000100000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000; // D (0x00000020000000000400000000000000) 
14'h12cb : LOC =         127'b0000000000000000000000001000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000; // D (0x00000040000000000400000000000000) 
14'h1f73 : LOC =         127'b0000000000000000000000010000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000; // D (0x00000080000000000400000000000000) 
14'h0403 : LOC =         127'b0000000000000000000000100000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000; // D (0x00000100000000000400000000000000) 
14'h32e3 : LOC =         127'b0000000000000000000001000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000; // D (0x00000200000000000400000000000000) 
14'h1c54 : LOC =         127'b0000000000000000000010000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000; // D (0x00000400000000000400000000000000) 
14'h024d : LOC =         127'b0000000000000000000100000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000; // D (0x00000800000000000400000000000000) 
14'h3e7f : LOC =         127'b0000000000000000001000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000; // D (0x00001000000000000400000000000000) 
14'h056c : LOC =         127'b0000000000000000010000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000; // D (0x00002000000000000400000000000000) 
14'h303d : LOC =         127'b0000000000000000100000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000; // D (0x00004000000000000400000000000000) 
14'h19e8 : LOC =         127'b0000000000000001000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000; // D (0x00008000000000000400000000000000) 
14'h0935 : LOC =         127'b0000000000000010000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000; // D (0x00010000000000000400000000000000) 
14'h288f : LOC =         127'b0000000000000100000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000; // D (0x00020000000000000400000000000000) 
14'h288c : LOC =         127'b0000000000001000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000; // D (0x00040000000000000400000000000000) 
14'h288a : LOC =         127'b0000000000010000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000; // D (0x00080000000000000400000000000000) 
14'h2886 : LOC =         127'b0000000000100000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000; // D (0x00100000000000000400000000000000) 
14'h289e : LOC =         127'b0000000001000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000; // D (0x00200000000000000400000000000000) 
14'h28ae : LOC =         127'b0000000010000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000; // D (0x00400000000000000400000000000000) 
14'h28ce : LOC =         127'b0000000100000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000; // D (0x00800000000000000400000000000000) 
14'h280e : LOC =         127'b0000001000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000; // D (0x01000000000000000400000000000000) 
14'h298e : LOC =         127'b0000010000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000; // D (0x02000000000000000400000000000000) 
14'h2a8e : LOC =         127'b0000100000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000; // D (0x04000000000000000400000000000000) 
14'h2c8e : LOC =         127'b0001000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000; // D (0x08000000000000000400000000000000) 
14'h208e : LOC =         127'b0010000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000; // D (0x10000000000000000400000000000000) 
14'h388e : LOC =         127'b0100000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000; // D (0x20000000000000000400000000000000) 
14'h088e : LOC =         127'b1000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000; // D (0x40000000000000000400000000000000) 
14'h126b : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000; // S (0x00000000000000000800000000000000) 
14'h36bd : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000; // D (0x00000000000000001800000000000000) 
14'h18b0 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000000000000000000000000000000000000; // D (0x00000000000000002800000000000000) 
14'h07dd : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000; // D (0x00000000000000004800000000000000) 
14'h3907 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000001000100000000000000000000000000000000000000000000000000000000000; // D (0x00000000000000008800000000000000) 
14'h07c4 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000010000100000000000000000000000000000000000000000000000000000000000; // D (0x00000000000000010800000000000000) 
14'h3935 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000100000100000000000000000000000000000000000000000000000000000000000; // D (0x00000000000000020800000000000000) 
14'h07a0 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000001000000100000000000000000000000000000000000000000000000000000000000; // D (0x00000000000000040800000000000000) 
14'h39fd : LOC =         127'b0000000000000000000000000000000000000000000000000000000000010000000100000000000000000000000000000000000000000000000000000000000; // D (0x00000000000000080800000000000000) 
14'h0630 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000100000000100000000000000000000000000000000000000000000000000000000000; // D (0x00000000000000100800000000000000) 
14'h3add : LOC =         127'b0000000000000000000000000000000000000000000000000000000001000000000100000000000000000000000000000000000000000000000000000000000; // D (0x00000000000000200800000000000000) 
14'h0070 : LOC =         127'b0000000000000000000000000000000000000000000000000000000010000000000100000000000000000000000000000000000000000000000000000000000; // D (0x00000000000000400800000000000000) 
14'h365d : LOC =         127'b0000000000000000000000000000000000000000000000000000000100000000000100000000000000000000000000000000000000000000000000000000000; // D (0x00000000000000800800000000000000) 
14'h1970 : LOC =         127'b0000000000000000000000000000000000000000000000000000001000000000000100000000000000000000000000000000000000000000000000000000000; // D (0x00000000000001000800000000000000) 
14'h045d : LOC =         127'b0000000000000000000000000000000000000000000000000000010000000000000100000000000000000000000000000000000000000000000000000000000; // D (0x00000000000002000800000000000000) 
14'h3e07 : LOC =         127'b0000000000000000000000000000000000000000000000000000100000000000000100000000000000000000000000000000000000000000000000000000000; // D (0x00000000000004000800000000000000) 
14'h09c4 : LOC =         127'b0000000000000000000000000000000000000000000000000001000000000000000100000000000000000000000000000000000000000000000000000000000; // D (0x00000000000008000800000000000000) 
14'h2535 : LOC =         127'b0000000000000000000000000000000000000000000000000010000000000000000100000000000000000000000000000000000000000000000000000000000; // D (0x00000000000010000800000000000000) 
14'h3fa0 : LOC =         127'b0000000000000000000000000000000000000000000000000100000000000000000100000000000000000000000000000000000000000000000000000000000; // D (0x00000000000020000800000000000000) 
14'h0a8a : LOC =         127'b0000000000000000000000000000000000000000000000001000000000000000000100000000000000000000000000000000000000000000000000000000000; // D (0x00000000000040000800000000000000) 
14'h23a9 : LOC =         127'b0000000000000000000000000000000000000000000000010000000000000000000100000000000000000000000000000000000000000000000000000000000; // D (0x00000000000080000800000000000000) 
14'h3298 : LOC =         127'b0000000000000000000000000000000000000000000000100000000000000000000100000000000000000000000000000000000000000000000000000000000; // D (0x00000000000100000800000000000000) 
14'h10fa : LOC =         127'b0000000000000000000000000000000000000000000001000000000000000000000100000000000000000000000000000000000000000000000000000000000; // D (0x00000000000200000800000000000000) 
14'h1749 : LOC =         127'b0000000000000000000000000000000000000000000010000000000000000000000100000000000000000000000000000000000000000000000000000000000; // D (0x00000000000400000800000000000000) 
14'h182f : LOC =         127'b0000000000000000000000000000000000000000000100000000000000000000000100000000000000000000000000000000000000000000000000000000000; // D (0x00000000000800000800000000000000) 
14'h06e3 : LOC =         127'b0000000000000000000000000000000000000000001000000000000000000000000100000000000000000000000000000000000000000000000000000000000; // D (0x00000000001000000800000000000000) 
14'h3b7b : LOC =         127'b0000000000000000000000000000000000000000010000000000000000000000000100000000000000000000000000000000000000000000000000000000000; // D (0x00000000002000000800000000000000) 
14'h033c : LOC =         127'b0000000000000000000000000000000000000000100000000000000000000000000100000000000000000000000000000000000000000000000000000000000; // D (0x00000000004000000800000000000000) 
14'h30c5 : LOC =         127'b0000000000000000000000000000000000000001000000000000000000000000000100000000000000000000000000000000000000000000000000000000000; // D (0x00000000008000000800000000000000) 
14'h1440 : LOC =         127'b0000000000000000000000000000000000000010000000000000000000000000000100000000000000000000000000000000000000000000000000000000000; // D (0x00000000010000000800000000000000) 
14'h1e3d : LOC =         127'b0000000000000000000000000000000000000100000000000000000000000000000100000000000000000000000000000000000000000000000000000000000; // D (0x00000000020000000800000000000000) 
14'h0ac7 : LOC =         127'b0000000000000000000000000000000000001000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000; // D (0x00000000040000000800000000000000) 
14'h2333 : LOC =         127'b0000000000000000000000000000000000010000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000; // D (0x00000000080000000800000000000000) 
14'h33ac : LOC =         127'b0000000000000000000000000000000000100000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000; // D (0x00000000100000000800000000000000) 
14'h1292 : LOC =         127'b0000000000000000000000000000000001000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000; // D (0x00000000200000000800000000000000) 
14'h1399 : LOC =         127'b0000000000000000000000000000000010000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000; // D (0x00000000400000000800000000000000) 
14'h118f : LOC =         127'b0000000000000000000000000000000100000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000; // D (0x00000000800000000800000000000000) 
14'h15a3 : LOC =         127'b0000000000000000000000000000001000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000; // D (0x00000001000000000800000000000000) 
14'h1dfb : LOC =         127'b0000000000000000000000000000010000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000; // D (0x00000002000000000800000000000000) 
14'h0d4b : LOC =         127'b0000000000000000000000000000100000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000; // D (0x00000004000000000800000000000000) 
14'h2c2b : LOC =         127'b0000000000000000000000000001000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000; // D (0x00000008000000000800000000000000) 
14'h2d9c : LOC =         127'b0000000000000000000000000010000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000; // D (0x00000010000000000800000000000000) 
14'h2ef2 : LOC =         127'b0000000000000000000000000100000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000; // D (0x00000020000000000800000000000000) 
14'h282e : LOC =         127'b0000000000000000000000001000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000; // D (0x00000040000000000800000000000000) 
14'h2596 : LOC =         127'b0000000000000000000000010000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000; // D (0x00000080000000000800000000000000) 
14'h3ee6 : LOC =         127'b0000000000000000000000100000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000; // D (0x00000100000000000800000000000000) 
14'h0806 : LOC =         127'b0000000000000000000001000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000; // D (0x00000200000000000800000000000000) 
14'h26b1 : LOC =         127'b0000000000000000000010000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000; // D (0x00000400000000000800000000000000) 
14'h38a8 : LOC =         127'b0000000000000000000100000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000; // D (0x00000800000000000800000000000000) 
14'h049a : LOC =         127'b0000000000000000001000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000; // D (0x00001000000000000800000000000000) 
14'h3f89 : LOC =         127'b0000000000000000010000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000; // D (0x00002000000000000800000000000000) 
14'h0ad8 : LOC =         127'b0000000000000000100000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000; // D (0x00004000000000000800000000000000) 
14'h230d : LOC =         127'b0000000000000001000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000; // D (0x00008000000000000800000000000000) 
14'h33d0 : LOC =         127'b0000000000000010000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000; // D (0x00010000000000000800000000000000) 
14'h126a : LOC =         127'b0000000000000100000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000; // D (0x00020000000000000800000000000000) 
14'h1269 : LOC =         127'b0000000000001000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000; // D (0x00040000000000000800000000000000) 
14'h126f : LOC =         127'b0000000000010000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000; // D (0x00080000000000000800000000000000) 
14'h1263 : LOC =         127'b0000000000100000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000; // D (0x00100000000000000800000000000000) 
14'h127b : LOC =         127'b0000000001000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000; // D (0x00200000000000000800000000000000) 
14'h124b : LOC =         127'b0000000010000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000; // D (0x00400000000000000800000000000000) 
14'h122b : LOC =         127'b0000000100000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000; // D (0x00800000000000000800000000000000) 
14'h12eb : LOC =         127'b0000001000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000; // D (0x01000000000000000800000000000000) 
14'h136b : LOC =         127'b0000010000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000; // D (0x02000000000000000800000000000000) 
14'h106b : LOC =         127'b0000100000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000; // D (0x04000000000000000800000000000000) 
14'h166b : LOC =         127'b0001000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000; // D (0x08000000000000000800000000000000) 
14'h1a6b : LOC =         127'b0010000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000; // D (0x10000000000000000800000000000000) 
14'h026b : LOC =         127'b0100000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000; // D (0x20000000000000000800000000000000) 
14'h326b : LOC =         127'b1000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000; // D (0x40000000000000000800000000000000) 
14'h24d6 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000; // S (0x00000000000000001000000000000000) 
14'h2e0d : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000000003000000000000000) 
14'h3160 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000101000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000000005000000000000000) 
14'h0fba : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000000009000000000000000) 
14'h3179 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000010001000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000000011000000000000000) 
14'h0f88 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000100001000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000000021000000000000000) 
14'h311d : LOC =         127'b0000000000000000000000000000000000000000000000000000000000001000001000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000000041000000000000000) 
14'h0f40 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000010000001000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000000081000000000000000) 
14'h308d : LOC =         127'b0000000000000000000000000000000000000000000000000000000000100000001000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000000101000000000000000) 
14'h0c60 : LOC =         127'b0000000000000000000000000000000000000000000000000000000001000000001000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000000201000000000000000) 
14'h36cd : LOC =         127'b0000000000000000000000000000000000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000000401000000000000000) 
14'h00e0 : LOC =         127'b0000000000000000000000000000000000000000000000000000000100000000001000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000000801000000000000000) 
14'h2fcd : LOC =         127'b0000000000000000000000000000000000000000000000000000001000000000001000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000001001000000000000000) 
14'h32e0 : LOC =         127'b0000000000000000000000000000000000000000000000000000010000000000001000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000002001000000000000000) 
14'h08ba : LOC =         127'b0000000000000000000000000000000000000000000000000000100000000000001000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000004001000000000000000) 
14'h3f79 : LOC =         127'b0000000000000000000000000000000000000000000000000001000000000000001000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000008001000000000000000) 
14'h1388 : LOC =         127'b0000000000000000000000000000000000000000000000000010000000000000001000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000010001000000000000000) 
14'h091d : LOC =         127'b0000000000000000000000000000000000000000000000000100000000000000001000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000020001000000000000000) 
14'h3c37 : LOC =         127'b0000000000000000000000000000000000000000000000001000000000000000001000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000040001000000000000000) 
14'h1514 : LOC =         127'b0000000000000000000000000000000000000000000000010000000000000000001000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000080001000000000000000) 
14'h0425 : LOC =         127'b0000000000000000000000000000000000000000000000100000000000000000001000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000100001000000000000000) 
14'h2647 : LOC =         127'b0000000000000000000000000000000000000000000001000000000000000000001000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000200001000000000000000) 
14'h21f4 : LOC =         127'b0000000000000000000000000000000000000000000010000000000000000000001000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000400001000000000000000) 
14'h2e92 : LOC =         127'b0000000000000000000000000000000000000000000100000000000000000000001000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000800001000000000000000) 
14'h305e : LOC =         127'b0000000000000000000000000000000000000000001000000000000000000000001000000000000000000000000000000000000000000000000000000000000; // D (0x00000000001000001000000000000000) 
14'h0dc6 : LOC =         127'b0000000000000000000000000000000000000000010000000000000000000000001000000000000000000000000000000000000000000000000000000000000; // D (0x00000000002000001000000000000000) 
14'h3581 : LOC =         127'b0000000000000000000000000000000000000000100000000000000000000000001000000000000000000000000000000000000000000000000000000000000; // D (0x00000000004000001000000000000000) 
14'h0678 : LOC =         127'b0000000000000000000000000000000000000001000000000000000000000000001000000000000000000000000000000000000000000000000000000000000; // D (0x00000000008000001000000000000000) 
14'h22fd : LOC =         127'b0000000000000000000000000000000000000010000000000000000000000000001000000000000000000000000000000000000000000000000000000000000; // D (0x00000000010000001000000000000000) 
14'h2880 : LOC =         127'b0000000000000000000000000000000000000100000000000000000000000000001000000000000000000000000000000000000000000000000000000000000; // D (0x00000000020000001000000000000000) 
14'h3c7a : LOC =         127'b0000000000000000000000000000000000001000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000; // D (0x00000000040000001000000000000000) 
14'h158e : LOC =         127'b0000000000000000000000000000000000010000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000; // D (0x00000000080000001000000000000000) 
14'h0511 : LOC =         127'b0000000000000000000000000000000000100000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000; // D (0x00000000100000001000000000000000) 
14'h242f : LOC =         127'b0000000000000000000000000000000001000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000; // D (0x00000000200000001000000000000000) 
14'h2524 : LOC =         127'b0000000000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000; // D (0x00000000400000001000000000000000) 
14'h2732 : LOC =         127'b0000000000000000000000000000000100000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000; // D (0x00000000800000001000000000000000) 
14'h231e : LOC =         127'b0000000000000000000000000000001000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000; // D (0x00000001000000001000000000000000) 
14'h2b46 : LOC =         127'b0000000000000000000000000000010000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000; // D (0x00000002000000001000000000000000) 
14'h3bf6 : LOC =         127'b0000000000000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000; // D (0x00000004000000001000000000000000) 
14'h1a96 : LOC =         127'b0000000000000000000000000001000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000; // D (0x00000008000000001000000000000000) 
14'h1b21 : LOC =         127'b0000000000000000000000000010000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000; // D (0x00000010000000001000000000000000) 
14'h184f : LOC =         127'b0000000000000000000000000100000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000; // D (0x00000020000000001000000000000000) 
14'h1e93 : LOC =         127'b0000000000000000000000001000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000; // D (0x00000040000000001000000000000000) 
14'h132b : LOC =         127'b0000000000000000000000010000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000; // D (0x00000080000000001000000000000000) 
14'h085b : LOC =         127'b0000000000000000000000100000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000; // D (0x00000100000000001000000000000000) 
14'h3ebb : LOC =         127'b0000000000000000000001000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000; // D (0x00000200000000001000000000000000) 
14'h100c : LOC =         127'b0000000000000000000010000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000; // D (0x00000400000000001000000000000000) 
14'h0e15 : LOC =         127'b0000000000000000000100000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000; // D (0x00000800000000001000000000000000) 
14'h3227 : LOC =         127'b0000000000000000001000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000; // D (0x00001000000000001000000000000000) 
14'h0934 : LOC =         127'b0000000000000000010000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000; // D (0x00002000000000001000000000000000) 
14'h3c65 : LOC =         127'b0000000000000000100000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000; // D (0x00004000000000001000000000000000) 
14'h15b0 : LOC =         127'b0000000000000001000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000; // D (0x00008000000000001000000000000000) 
14'h056d : LOC =         127'b0000000000000010000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000; // D (0x00010000000000001000000000000000) 
14'h24d7 : LOC =         127'b0000000000000100000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000; // D (0x00020000000000001000000000000000) 
14'h24d4 : LOC =         127'b0000000000001000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000; // D (0x00040000000000001000000000000000) 
14'h24d2 : LOC =         127'b0000000000010000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000; // D (0x00080000000000001000000000000000) 
14'h24de : LOC =         127'b0000000000100000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000; // D (0x00100000000000001000000000000000) 
14'h24c6 : LOC =         127'b0000000001000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000; // D (0x00200000000000001000000000000000) 
14'h24f6 : LOC =         127'b0000000010000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000; // D (0x00400000000000001000000000000000) 
14'h2496 : LOC =         127'b0000000100000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000; // D (0x00800000000000001000000000000000) 
14'h2456 : LOC =         127'b0000001000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000; // D (0x01000000000000001000000000000000) 
14'h25d6 : LOC =         127'b0000010000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000; // D (0x02000000000000001000000000000000) 
14'h26d6 : LOC =         127'b0000100000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000; // D (0x04000000000000001000000000000000) 
14'h20d6 : LOC =         127'b0001000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000; // D (0x08000000000000001000000000000000) 
14'h2cd6 : LOC =         127'b0010000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000; // D (0x10000000000000001000000000000000) 
14'h34d6 : LOC =         127'b0100000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000; // D (0x20000000000000001000000000000000) 
14'h04d6 : LOC =         127'b1000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000; // D (0x40000000000000001000000000000000) 
14'h0adb : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000; // S (0x00000000000000002000000000000000) 
14'h1f6d : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000000006000000000000000) 
14'h21b7 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000001010000000000000000000000000000000000000000000000000000000000000; // D (0x0000000000000000a000000000000000) 
14'h1f74 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000000012000000000000000) 
14'h2185 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000100010000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000000022000000000000000) 
14'h1f10 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000001000010000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000000042000000000000000) 
14'h214d : LOC =         127'b0000000000000000000000000000000000000000000000000000000000010000010000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000000082000000000000000) 
14'h1e80 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000100000010000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000000102000000000000000) 
14'h226d : LOC =         127'b0000000000000000000000000000000000000000000000000000000001000000010000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000000202000000000000000) 
14'h18c0 : LOC =         127'b0000000000000000000000000000000000000000000000000000000010000000010000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000000402000000000000000) 
14'h2eed : LOC =         127'b0000000000000000000000000000000000000000000000000000000100000000010000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000000802000000000000000) 
14'h01c0 : LOC =         127'b0000000000000000000000000000000000000000000000000000001000000000010000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000001002000000000000000) 
14'h1ced : LOC =         127'b0000000000000000000000000000000000000000000000000000010000000000010000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000002002000000000000000) 
14'h26b7 : LOC =         127'b0000000000000000000000000000000000000000000000000000100000000000010000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000004002000000000000000) 
14'h1174 : LOC =         127'b0000000000000000000000000000000000000000000000000001000000000000010000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000008002000000000000000) 
14'h3d85 : LOC =         127'b0000000000000000000000000000000000000000000000000010000000000000010000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000010002000000000000000) 
14'h2710 : LOC =         127'b0000000000000000000000000000000000000000000000000100000000000000010000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000020002000000000000000) 
14'h123a : LOC =         127'b0000000000000000000000000000000000000000000000001000000000000000010000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000040002000000000000000) 
14'h3b19 : LOC =         127'b0000000000000000000000000000000000000000000000010000000000000000010000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000080002000000000000000) 
14'h2a28 : LOC =         127'b0000000000000000000000000000000000000000000000100000000000000000010000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000100002000000000000000) 
14'h084a : LOC =         127'b0000000000000000000000000000000000000000000001000000000000000000010000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000200002000000000000000) 
14'h0ff9 : LOC =         127'b0000000000000000000000000000000000000000000010000000000000000000010000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000400002000000000000000) 
14'h009f : LOC =         127'b0000000000000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000800002000000000000000) 
14'h1e53 : LOC =         127'b0000000000000000000000000000000000000000001000000000000000000000010000000000000000000000000000000000000000000000000000000000000; // D (0x00000000001000002000000000000000) 
14'h23cb : LOC =         127'b0000000000000000000000000000000000000000010000000000000000000000010000000000000000000000000000000000000000000000000000000000000; // D (0x00000000002000002000000000000000) 
14'h1b8c : LOC =         127'b0000000000000000000000000000000000000000100000000000000000000000010000000000000000000000000000000000000000000000000000000000000; // D (0x00000000004000002000000000000000) 
14'h2875 : LOC =         127'b0000000000000000000000000000000000000001000000000000000000000000010000000000000000000000000000000000000000000000000000000000000; // D (0x00000000008000002000000000000000) 
14'h0cf0 : LOC =         127'b0000000000000000000000000000000000000010000000000000000000000000010000000000000000000000000000000000000000000000000000000000000; // D (0x00000000010000002000000000000000) 
14'h068d : LOC =         127'b0000000000000000000000000000000000000100000000000000000000000000010000000000000000000000000000000000000000000000000000000000000; // D (0x00000000020000002000000000000000) 
14'h1277 : LOC =         127'b0000000000000000000000000000000000001000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000; // D (0x00000000040000002000000000000000) 
14'h3b83 : LOC =         127'b0000000000000000000000000000000000010000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000; // D (0x00000000080000002000000000000000) 
14'h2b1c : LOC =         127'b0000000000000000000000000000000000100000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000; // D (0x00000000100000002000000000000000) 
14'h0a22 : LOC =         127'b0000000000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000; // D (0x00000000200000002000000000000000) 
14'h0b29 : LOC =         127'b0000000000000000000000000000000010000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000; // D (0x00000000400000002000000000000000) 
14'h093f : LOC =         127'b0000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000; // D (0x00000000800000002000000000000000) 
14'h0d13 : LOC =         127'b0000000000000000000000000000001000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000; // D (0x00000001000000002000000000000000) 
14'h054b : LOC =         127'b0000000000000000000000000000010000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000; // D (0x00000002000000002000000000000000) 
14'h15fb : LOC =         127'b0000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000; // D (0x00000004000000002000000000000000) 
14'h349b : LOC =         127'b0000000000000000000000000001000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000; // D (0x00000008000000002000000000000000) 
14'h352c : LOC =         127'b0000000000000000000000000010000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000; // D (0x00000010000000002000000000000000) 
14'h3642 : LOC =         127'b0000000000000000000000000100000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000; // D (0x00000020000000002000000000000000) 
14'h309e : LOC =         127'b0000000000000000000000001000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000; // D (0x00000040000000002000000000000000) 
14'h3d26 : LOC =         127'b0000000000000000000000010000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000; // D (0x00000080000000002000000000000000) 
14'h2656 : LOC =         127'b0000000000000000000000100000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000; // D (0x00000100000000002000000000000000) 
14'h10b6 : LOC =         127'b0000000000000000000001000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000; // D (0x00000200000000002000000000000000) 
14'h3e01 : LOC =         127'b0000000000000000000010000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000; // D (0x00000400000000002000000000000000) 
14'h2018 : LOC =         127'b0000000000000000000100000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000; // D (0x00000800000000002000000000000000) 
14'h1c2a : LOC =         127'b0000000000000000001000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000; // D (0x00001000000000002000000000000000) 
14'h2739 : LOC =         127'b0000000000000000010000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000; // D (0x00002000000000002000000000000000) 
14'h1268 : LOC =         127'b0000000000000000100000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000; // D (0x00004000000000002000000000000000) 
14'h3bbd : LOC =         127'b0000000000000001000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000; // D (0x00008000000000002000000000000000) 
14'h2b60 : LOC =         127'b0000000000000010000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000; // D (0x00010000000000002000000000000000) 
14'h0ada : LOC =         127'b0000000000000100000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000; // D (0x00020000000000002000000000000000) 
14'h0ad9 : LOC =         127'b0000000000001000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000; // D (0x00040000000000002000000000000000) 
14'h0adf : LOC =         127'b0000000000010000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000; // D (0x00080000000000002000000000000000) 
14'h0ad3 : LOC =         127'b0000000000100000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000; // D (0x00100000000000002000000000000000) 
14'h0acb : LOC =         127'b0000000001000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000; // D (0x00200000000000002000000000000000) 
14'h0afb : LOC =         127'b0000000010000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000; // D (0x00400000000000002000000000000000) 
14'h0a9b : LOC =         127'b0000000100000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000; // D (0x00800000000000002000000000000000) 
14'h0a5b : LOC =         127'b0000001000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000; // D (0x01000000000000002000000000000000) 
14'h0bdb : LOC =         127'b0000010000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000; // D (0x02000000000000002000000000000000) 
14'h08db : LOC =         127'b0000100000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000; // D (0x04000000000000002000000000000000) 
14'h0edb : LOC =         127'b0001000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000; // D (0x08000000000000002000000000000000) 
14'h02db : LOC =         127'b0010000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000; // D (0x10000000000000002000000000000000) 
14'h1adb : LOC =         127'b0100000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000; // D (0x20000000000000002000000000000000) 
14'h2adb : LOC =         127'b1000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000; // D (0x40000000000000002000000000000000) 
14'h15b6 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000; // S (0x00000000000000004000000000000000) 
14'h3eda : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000; // D (0x0000000000000000c000000000000000) 
14'h0019 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000000014000000000000000) 
14'h3ee8 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000000024000000000000000) 
14'h007d : LOC =         127'b0000000000000000000000000000000000000000000000000000000000001000100000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000000044000000000000000) 
14'h3e20 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000010000100000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000000084000000000000000) 
14'h01ed : LOC =         127'b0000000000000000000000000000000000000000000000000000000000100000100000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000000104000000000000000) 
14'h3d00 : LOC =         127'b0000000000000000000000000000000000000000000000000000000001000000100000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000000204000000000000000) 
14'h07ad : LOC =         127'b0000000000000000000000000000000000000000000000000000000010000000100000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000000404000000000000000) 
14'h3180 : LOC =         127'b0000000000000000000000000000000000000000000000000000000100000000100000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000000804000000000000000) 
14'h1ead : LOC =         127'b0000000000000000000000000000000000000000000000000000001000000000100000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000001004000000000000000) 
14'h0380 : LOC =         127'b0000000000000000000000000000000000000000000000000000010000000000100000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000002004000000000000000) 
14'h39da : LOC =         127'b0000000000000000000000000000000000000000000000000000100000000000100000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000004004000000000000000) 
14'h0e19 : LOC =         127'b0000000000000000000000000000000000000000000000000001000000000000100000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000008004000000000000000) 
14'h22e8 : LOC =         127'b0000000000000000000000000000000000000000000000000010000000000000100000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000010004000000000000000) 
14'h387d : LOC =         127'b0000000000000000000000000000000000000000000000000100000000000000100000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000020004000000000000000) 
14'h0d57 : LOC =         127'b0000000000000000000000000000000000000000000000001000000000000000100000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000040004000000000000000) 
14'h2474 : LOC =         127'b0000000000000000000000000000000000000000000000010000000000000000100000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000080004000000000000000) 
14'h3545 : LOC =         127'b0000000000000000000000000000000000000000000000100000000000000000100000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000100004000000000000000) 
14'h1727 : LOC =         127'b0000000000000000000000000000000000000000000001000000000000000000100000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000200004000000000000000) 
14'h1094 : LOC =         127'b0000000000000000000000000000000000000000000010000000000000000000100000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000400004000000000000000) 
14'h1ff2 : LOC =         127'b0000000000000000000000000000000000000000000100000000000000000000100000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000800004000000000000000) 
14'h013e : LOC =         127'b0000000000000000000000000000000000000000001000000000000000000000100000000000000000000000000000000000000000000000000000000000000; // D (0x00000000001000004000000000000000) 
14'h3ca6 : LOC =         127'b0000000000000000000000000000000000000000010000000000000000000000100000000000000000000000000000000000000000000000000000000000000; // D (0x00000000002000004000000000000000) 
14'h04e1 : LOC =         127'b0000000000000000000000000000000000000000100000000000000000000000100000000000000000000000000000000000000000000000000000000000000; // D (0x00000000004000004000000000000000) 
14'h3718 : LOC =         127'b0000000000000000000000000000000000000001000000000000000000000000100000000000000000000000000000000000000000000000000000000000000; // D (0x00000000008000004000000000000000) 
14'h139d : LOC =         127'b0000000000000000000000000000000000000010000000000000000000000000100000000000000000000000000000000000000000000000000000000000000; // D (0x00000000010000004000000000000000) 
14'h19e0 : LOC =         127'b0000000000000000000000000000000000000100000000000000000000000000100000000000000000000000000000000000000000000000000000000000000; // D (0x00000000020000004000000000000000) 
14'h0d1a : LOC =         127'b0000000000000000000000000000000000001000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000; // D (0x00000000040000004000000000000000) 
14'h24ee : LOC =         127'b0000000000000000000000000000000000010000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000; // D (0x00000000080000004000000000000000) 
14'h3471 : LOC =         127'b0000000000000000000000000000000000100000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000; // D (0x00000000100000004000000000000000) 
14'h154f : LOC =         127'b0000000000000000000000000000000001000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000; // D (0x00000000200000004000000000000000) 
14'h1444 : LOC =         127'b0000000000000000000000000000000010000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000; // D (0x00000000400000004000000000000000) 
14'h1652 : LOC =         127'b0000000000000000000000000000000100000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000; // D (0x00000000800000004000000000000000) 
14'h127e : LOC =         127'b0000000000000000000000000000001000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000; // D (0x00000001000000004000000000000000) 
14'h1a26 : LOC =         127'b0000000000000000000000000000010000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000; // D (0x00000002000000004000000000000000) 
14'h0a96 : LOC =         127'b0000000000000000000000000000100000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000; // D (0x00000004000000004000000000000000) 
14'h2bf6 : LOC =         127'b0000000000000000000000000001000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000; // D (0x00000008000000004000000000000000) 
14'h2a41 : LOC =         127'b0000000000000000000000000010000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000; // D (0x00000010000000004000000000000000) 
14'h292f : LOC =         127'b0000000000000000000000000100000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000; // D (0x00000020000000004000000000000000) 
14'h2ff3 : LOC =         127'b0000000000000000000000001000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000; // D (0x00000040000000004000000000000000) 
14'h224b : LOC =         127'b0000000000000000000000010000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000; // D (0x00000080000000004000000000000000) 
14'h393b : LOC =         127'b0000000000000000000000100000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000; // D (0x00000100000000004000000000000000) 
14'h0fdb : LOC =         127'b0000000000000000000001000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000; // D (0x00000200000000004000000000000000) 
14'h216c : LOC =         127'b0000000000000000000010000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000; // D (0x00000400000000004000000000000000) 
14'h3f75 : LOC =         127'b0000000000000000000100000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000; // D (0x00000800000000004000000000000000) 
14'h0347 : LOC =         127'b0000000000000000001000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000; // D (0x00001000000000004000000000000000) 
14'h3854 : LOC =         127'b0000000000000000010000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000; // D (0x00002000000000004000000000000000) 
14'h0d05 : LOC =         127'b0000000000000000100000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000; // D (0x00004000000000004000000000000000) 
14'h24d0 : LOC =         127'b0000000000000001000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000; // D (0x00008000000000004000000000000000) 
14'h340d : LOC =         127'b0000000000000010000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000; // D (0x00010000000000004000000000000000) 
14'h15b7 : LOC =         127'b0000000000000100000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000; // D (0x00020000000000004000000000000000) 
14'h15b4 : LOC =         127'b0000000000001000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000; // D (0x00040000000000004000000000000000) 
14'h15b2 : LOC =         127'b0000000000010000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000; // D (0x00080000000000004000000000000000) 
14'h15be : LOC =         127'b0000000000100000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000; // D (0x00100000000000004000000000000000) 
14'h15a6 : LOC =         127'b0000000001000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000; // D (0x00200000000000004000000000000000) 
14'h1596 : LOC =         127'b0000000010000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000; // D (0x00400000000000004000000000000000) 
14'h15f6 : LOC =         127'b0000000100000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000; // D (0x00800000000000004000000000000000) 
14'h1536 : LOC =         127'b0000001000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000; // D (0x01000000000000004000000000000000) 
14'h14b6 : LOC =         127'b0000010000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000; // D (0x02000000000000004000000000000000) 
14'h17b6 : LOC =         127'b0000100000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000; // D (0x04000000000000004000000000000000) 
14'h11b6 : LOC =         127'b0001000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000; // D (0x08000000000000004000000000000000) 
14'h1db6 : LOC =         127'b0010000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000; // D (0x10000000000000004000000000000000) 
14'h05b6 : LOC =         127'b0100000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000; // D (0x20000000000000004000000000000000) 
14'h35b6 : LOC =         127'b1000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000; // D (0x40000000000000004000000000000000) 
14'h2b6c : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000; // S (0x00000000000000008000000000000000) 
14'h3ec3 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000011000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000000018000000000000000) 
14'h0032 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000101000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000000028000000000000000) 
14'h3ea7 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000000048000000000000000) 
14'h00fa : LOC =         127'b0000000000000000000000000000000000000000000000000000000000010001000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000000088000000000000000) 
14'h3f37 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000100001000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000000108000000000000000) 
14'h03da : LOC =         127'b0000000000000000000000000000000000000000000000000000000001000001000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000000208000000000000000) 
14'h3977 : LOC =         127'b0000000000000000000000000000000000000000000000000000000010000001000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000000408000000000000000) 
14'h0f5a : LOC =         127'b0000000000000000000000000000000000000000000000000000000100000001000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000000808000000000000000) 
14'h2077 : LOC =         127'b0000000000000000000000000000000000000000000000000000001000000001000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000001008000000000000000) 
14'h3d5a : LOC =         127'b0000000000000000000000000000000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000002008000000000000000) 
14'h0700 : LOC =         127'b0000000000000000000000000000000000000000000000000000100000000001000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000004008000000000000000) 
14'h30c3 : LOC =         127'b0000000000000000000000000000000000000000000000000001000000000001000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000008008000000000000000) 
14'h1c32 : LOC =         127'b0000000000000000000000000000000000000000000000000010000000000001000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000010008000000000000000) 
14'h06a7 : LOC =         127'b0000000000000000000000000000000000000000000000000100000000000001000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000020008000000000000000) 
14'h338d : LOC =         127'b0000000000000000000000000000000000000000000000001000000000000001000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000040008000000000000000) 
14'h1aae : LOC =         127'b0000000000000000000000000000000000000000000000010000000000000001000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000080008000000000000000) 
14'h0b9f : LOC =         127'b0000000000000000000000000000000000000000000000100000000000000001000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000100008000000000000000) 
14'h29fd : LOC =         127'b0000000000000000000000000000000000000000000001000000000000000001000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000200008000000000000000) 
14'h2e4e : LOC =         127'b0000000000000000000000000000000000000000000010000000000000000001000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000400008000000000000000) 
14'h2128 : LOC =         127'b0000000000000000000000000000000000000000000100000000000000000001000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000800008000000000000000) 
14'h3fe4 : LOC =         127'b0000000000000000000000000000000000000000001000000000000000000001000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000001000008000000000000000) 
14'h027c : LOC =         127'b0000000000000000000000000000000000000000010000000000000000000001000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000002000008000000000000000) 
14'h3a3b : LOC =         127'b0000000000000000000000000000000000000000100000000000000000000001000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000004000008000000000000000) 
14'h09c2 : LOC =         127'b0000000000000000000000000000000000000001000000000000000000000001000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000008000008000000000000000) 
14'h2d47 : LOC =         127'b0000000000000000000000000000000000000010000000000000000000000001000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000010000008000000000000000) 
14'h273a : LOC =         127'b0000000000000000000000000000000000000100000000000000000000000001000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000020000008000000000000000) 
14'h33c0 : LOC =         127'b0000000000000000000000000000000000001000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000040000008000000000000000) 
14'h1a34 : LOC =         127'b0000000000000000000000000000000000010000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000080000008000000000000000) 
14'h0aab : LOC =         127'b0000000000000000000000000000000000100000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000100000008000000000000000) 
14'h2b95 : LOC =         127'b0000000000000000000000000000000001000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000200000008000000000000000) 
14'h2a9e : LOC =         127'b0000000000000000000000000000000010000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000400000008000000000000000) 
14'h2888 : LOC =         127'b0000000000000000000000000000000100000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000800000008000000000000000) 
14'h2ca4 : LOC =         127'b0000000000000000000000000000001000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000; // D (0x00000001000000008000000000000000) 
14'h24fc : LOC =         127'b0000000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000; // D (0x00000002000000008000000000000000) 
14'h344c : LOC =         127'b0000000000000000000000000000100000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000; // D (0x00000004000000008000000000000000) 
14'h152c : LOC =         127'b0000000000000000000000000001000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000; // D (0x00000008000000008000000000000000) 
14'h149b : LOC =         127'b0000000000000000000000000010000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000; // D (0x00000010000000008000000000000000) 
14'h17f5 : LOC =         127'b0000000000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000; // D (0x00000020000000008000000000000000) 
14'h1129 : LOC =         127'b0000000000000000000000001000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000; // D (0x00000040000000008000000000000000) 
14'h1c91 : LOC =         127'b0000000000000000000000010000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000; // D (0x00000080000000008000000000000000) 
14'h07e1 : LOC =         127'b0000000000000000000000100000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000; // D (0x00000100000000008000000000000000) 
14'h3101 : LOC =         127'b0000000000000000000001000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000; // D (0x00000200000000008000000000000000) 
14'h1fb6 : LOC =         127'b0000000000000000000010000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000; // D (0x00000400000000008000000000000000) 
14'h01af : LOC =         127'b0000000000000000000100000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000; // D (0x00000800000000008000000000000000) 
14'h3d9d : LOC =         127'b0000000000000000001000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000; // D (0x00001000000000008000000000000000) 
14'h068e : LOC =         127'b0000000000000000010000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000; // D (0x00002000000000008000000000000000) 
14'h33df : LOC =         127'b0000000000000000100000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000; // D (0x00004000000000008000000000000000) 
14'h1a0a : LOC =         127'b0000000000000001000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000; // D (0x00008000000000008000000000000000) 
14'h0ad7 : LOC =         127'b0000000000000010000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000; // D (0x00010000000000008000000000000000) 
14'h2b6d : LOC =         127'b0000000000000100000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000; // D (0x00020000000000008000000000000000) 
14'h2b6e : LOC =         127'b0000000000001000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000; // D (0x00040000000000008000000000000000) 
14'h2b68 : LOC =         127'b0000000000010000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000; // D (0x00080000000000008000000000000000) 
14'h2b64 : LOC =         127'b0000000000100000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000; // D (0x00100000000000008000000000000000) 
14'h2b7c : LOC =         127'b0000000001000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000; // D (0x00200000000000008000000000000000) 
14'h2b4c : LOC =         127'b0000000010000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000; // D (0x00400000000000008000000000000000) 
14'h2b2c : LOC =         127'b0000000100000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000; // D (0x00800000000000008000000000000000) 
14'h2bec : LOC =         127'b0000001000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000; // D (0x01000000000000008000000000000000) 
14'h2a6c : LOC =         127'b0000010000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000; // D (0x02000000000000008000000000000000) 
14'h296c : LOC =         127'b0000100000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000; // D (0x04000000000000008000000000000000) 
14'h2f6c : LOC =         127'b0001000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000; // D (0x08000000000000008000000000000000) 
14'h236c : LOC =         127'b0010000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000; // D (0x10000000000000008000000000000000) 
14'h3b6c : LOC =         127'b0100000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000; // D (0x20000000000000008000000000000000) 
14'h0b6c : LOC =         127'b1000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000; // D (0x40000000000000008000000000000000) 
14'h15af : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000; // S (0x00000000000000010000000000000000) 
14'h3ef1 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000000030000000000000000) 
14'h0064 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000001010000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000000050000000000000000) 
14'h3e39 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000000090000000000000000) 
14'h01f4 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000100010000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000000110000000000000000) 
14'h3d19 : LOC =         127'b0000000000000000000000000000000000000000000000000000000001000010000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000000210000000000000000) 
14'h07b4 : LOC =         127'b0000000000000000000000000000000000000000000000000000000010000010000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000000410000000000000000) 
14'h3199 : LOC =         127'b0000000000000000000000000000000000000000000000000000000100000010000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000000810000000000000000) 
14'h1eb4 : LOC =         127'b0000000000000000000000000000000000000000000000000000001000000010000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000001010000000000000000) 
14'h0399 : LOC =         127'b0000000000000000000000000000000000000000000000000000010000000010000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000002010000000000000000) 
14'h39c3 : LOC =         127'b0000000000000000000000000000000000000000000000000000100000000010000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000004010000000000000000) 
14'h0e00 : LOC =         127'b0000000000000000000000000000000000000000000000000001000000000010000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000008010000000000000000) 
14'h22f1 : LOC =         127'b0000000000000000000000000000000000000000000000000010000000000010000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000010010000000000000000) 
14'h3864 : LOC =         127'b0000000000000000000000000000000000000000000000000100000000000010000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000020010000000000000000) 
14'h0d4e : LOC =         127'b0000000000000000000000000000000000000000000000001000000000000010000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000040010000000000000000) 
14'h246d : LOC =         127'b0000000000000000000000000000000000000000000000010000000000000010000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000080010000000000000000) 
14'h355c : LOC =         127'b0000000000000000000000000000000000000000000000100000000000000010000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000100010000000000000000) 
14'h173e : LOC =         127'b0000000000000000000000000000000000000000000001000000000000000010000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000200010000000000000000) 
14'h108d : LOC =         127'b0000000000000000000000000000000000000000000010000000000000000010000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000400010000000000000000) 
14'h1feb : LOC =         127'b0000000000000000000000000000000000000000000100000000000000000010000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000800010000000000000000) 
14'h0127 : LOC =         127'b0000000000000000000000000000000000000000001000000000000000000010000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000001000010000000000000000) 
14'h3cbf : LOC =         127'b0000000000000000000000000000000000000000010000000000000000000010000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000002000010000000000000000) 
14'h04f8 : LOC =         127'b0000000000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000004000010000000000000000) 
14'h3701 : LOC =         127'b0000000000000000000000000000000000000001000000000000000000000010000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000008000010000000000000000) 
14'h1384 : LOC =         127'b0000000000000000000000000000000000000010000000000000000000000010000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000010000010000000000000000) 
14'h19f9 : LOC =         127'b0000000000000000000000000000000000000100000000000000000000000010000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000020000010000000000000000) 
14'h0d03 : LOC =         127'b0000000000000000000000000000000000001000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000040000010000000000000000) 
14'h24f7 : LOC =         127'b0000000000000000000000000000000000010000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000080000010000000000000000) 
14'h3468 : LOC =         127'b0000000000000000000000000000000000100000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000100000010000000000000000) 
14'h1556 : LOC =         127'b0000000000000000000000000000000001000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000200000010000000000000000) 
14'h145d : LOC =         127'b0000000000000000000000000000000010000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000400000010000000000000000) 
14'h164b : LOC =         127'b0000000000000000000000000000000100000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000800000010000000000000000) 
14'h1267 : LOC =         127'b0000000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000; // D (0x00000001000000010000000000000000) 
14'h1a3f : LOC =         127'b0000000000000000000000000000010000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000; // D (0x00000002000000010000000000000000) 
14'h0a8f : LOC =         127'b0000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000; // D (0x00000004000000010000000000000000) 
14'h2bef : LOC =         127'b0000000000000000000000000001000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000; // D (0x00000008000000010000000000000000) 
14'h2a58 : LOC =         127'b0000000000000000000000000010000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000; // D (0x00000010000000010000000000000000) 
14'h2936 : LOC =         127'b0000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000; // D (0x00000020000000010000000000000000) 
14'h2fea : LOC =         127'b0000000000000000000000001000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000; // D (0x00000040000000010000000000000000) 
14'h2252 : LOC =         127'b0000000000000000000000010000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000; // D (0x00000080000000010000000000000000) 
14'h3922 : LOC =         127'b0000000000000000000000100000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000; // D (0x00000100000000010000000000000000) 
14'h0fc2 : LOC =         127'b0000000000000000000001000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000; // D (0x00000200000000010000000000000000) 
14'h2175 : LOC =         127'b0000000000000000000010000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000; // D (0x00000400000000010000000000000000) 
14'h3f6c : LOC =         127'b0000000000000000000100000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000; // D (0x00000800000000010000000000000000) 
14'h035e : LOC =         127'b0000000000000000001000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000; // D (0x00001000000000010000000000000000) 
14'h384d : LOC =         127'b0000000000000000010000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000; // D (0x00002000000000010000000000000000) 
14'h0d1c : LOC =         127'b0000000000000000100000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000; // D (0x00004000000000010000000000000000) 
14'h24c9 : LOC =         127'b0000000000000001000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000; // D (0x00008000000000010000000000000000) 
14'h3414 : LOC =         127'b0000000000000010000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000; // D (0x00010000000000010000000000000000) 
14'h15ae : LOC =         127'b0000000000000100000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000; // D (0x00020000000000010000000000000000) 
14'h15ad : LOC =         127'b0000000000001000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000; // D (0x00040000000000010000000000000000) 
14'h15ab : LOC =         127'b0000000000010000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000; // D (0x00080000000000010000000000000000) 
14'h15a7 : LOC =         127'b0000000000100000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000; // D (0x00100000000000010000000000000000) 
14'h15bf : LOC =         127'b0000000001000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000; // D (0x00200000000000010000000000000000) 
14'h158f : LOC =         127'b0000000010000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000; // D (0x00400000000000010000000000000000) 
14'h15ef : LOC =         127'b0000000100000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000; // D (0x00800000000000010000000000000000) 
14'h152f : LOC =         127'b0000001000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000; // D (0x01000000000000010000000000000000) 
14'h14af : LOC =         127'b0000010000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000; // D (0x02000000000000010000000000000000) 
14'h17af : LOC =         127'b0000100000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000; // D (0x04000000000000010000000000000000) 
14'h11af : LOC =         127'b0001000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000; // D (0x08000000000000010000000000000000) 
14'h1daf : LOC =         127'b0010000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000; // D (0x10000000000000010000000000000000) 
14'h05af : LOC =         127'b0100000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000; // D (0x20000000000000010000000000000000) 
14'h35af : LOC =         127'b1000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000; // D (0x40000000000000010000000000000000) 
14'h2b5e : LOC =         127'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000; // S (0x00000000000000020000000000000000) 
14'h3e95 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000000060000000000000000) 
14'h00c8 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000010100000000000000000000000000000000000000000000000000000000000000000; // D (0x000000000000000a0000000000000000) 
14'h3f05 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000000120000000000000000) 
14'h03e8 : LOC =         127'b0000000000000000000000000000000000000000000000000000000001000100000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000000220000000000000000) 
14'h3945 : LOC =         127'b0000000000000000000000000000000000000000000000000000000010000100000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000000420000000000000000) 
14'h0f68 : LOC =         127'b0000000000000000000000000000000000000000000000000000000100000100000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000000820000000000000000) 
14'h2045 : LOC =         127'b0000000000000000000000000000000000000000000000000000001000000100000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000001020000000000000000) 
14'h3d68 : LOC =         127'b0000000000000000000000000000000000000000000000000000010000000100000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000002020000000000000000) 
14'h0732 : LOC =         127'b0000000000000000000000000000000000000000000000000000100000000100000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000004020000000000000000) 
14'h30f1 : LOC =         127'b0000000000000000000000000000000000000000000000000001000000000100000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000008020000000000000000) 
14'h1c00 : LOC =         127'b0000000000000000000000000000000000000000000000000010000000000100000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000010020000000000000000) 
14'h0695 : LOC =         127'b0000000000000000000000000000000000000000000000000100000000000100000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000020020000000000000000) 
14'h33bf : LOC =         127'b0000000000000000000000000000000000000000000000001000000000000100000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000040020000000000000000) 
14'h1a9c : LOC =         127'b0000000000000000000000000000000000000000000000010000000000000100000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000080020000000000000000) 
14'h0bad : LOC =         127'b0000000000000000000000000000000000000000000000100000000000000100000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000100020000000000000000) 
14'h29cf : LOC =         127'b0000000000000000000000000000000000000000000001000000000000000100000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000200020000000000000000) 
14'h2e7c : LOC =         127'b0000000000000000000000000000000000000000000010000000000000000100000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000400020000000000000000) 
14'h211a : LOC =         127'b0000000000000000000000000000000000000000000100000000000000000100000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000800020000000000000000) 
14'h3fd6 : LOC =         127'b0000000000000000000000000000000000000000001000000000000000000100000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000001000020000000000000000) 
14'h024e : LOC =         127'b0000000000000000000000000000000000000000010000000000000000000100000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000002000020000000000000000) 
14'h3a09 : LOC =         127'b0000000000000000000000000000000000000000100000000000000000000100000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000004000020000000000000000) 
14'h09f0 : LOC =         127'b0000000000000000000000000000000000000001000000000000000000000100000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000008000020000000000000000) 
14'h2d75 : LOC =         127'b0000000000000000000000000000000000000010000000000000000000000100000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000010000020000000000000000) 
14'h2708 : LOC =         127'b0000000000000000000000000000000000000100000000000000000000000100000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000020000020000000000000000) 
14'h33f2 : LOC =         127'b0000000000000000000000000000000000001000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000040000020000000000000000) 
14'h1a06 : LOC =         127'b0000000000000000000000000000000000010000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000080000020000000000000000) 
14'h0a99 : LOC =         127'b0000000000000000000000000000000000100000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000100000020000000000000000) 
14'h2ba7 : LOC =         127'b0000000000000000000000000000000001000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000200000020000000000000000) 
14'h2aac : LOC =         127'b0000000000000000000000000000000010000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000400000020000000000000000) 
14'h28ba : LOC =         127'b0000000000000000000000000000000100000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000800000020000000000000000) 
14'h2c96 : LOC =         127'b0000000000000000000000000000001000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000; // D (0x00000001000000020000000000000000) 
14'h24ce : LOC =         127'b0000000000000000000000000000010000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000; // D (0x00000002000000020000000000000000) 
14'h347e : LOC =         127'b0000000000000000000000000000100000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000; // D (0x00000004000000020000000000000000) 
14'h151e : LOC =         127'b0000000000000000000000000001000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000; // D (0x00000008000000020000000000000000) 
14'h14a9 : LOC =         127'b0000000000000000000000000010000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000; // D (0x00000010000000020000000000000000) 
14'h17c7 : LOC =         127'b0000000000000000000000000100000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000; // D (0x00000020000000020000000000000000) 
14'h111b : LOC =         127'b0000000000000000000000001000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000; // D (0x00000040000000020000000000000000) 
14'h1ca3 : LOC =         127'b0000000000000000000000010000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000; // D (0x00000080000000020000000000000000) 
14'h07d3 : LOC =         127'b0000000000000000000000100000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000; // D (0x00000100000000020000000000000000) 
14'h3133 : LOC =         127'b0000000000000000000001000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000; // D (0x00000200000000020000000000000000) 
14'h1f84 : LOC =         127'b0000000000000000000010000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000; // D (0x00000400000000020000000000000000) 
14'h019d : LOC =         127'b0000000000000000000100000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000; // D (0x00000800000000020000000000000000) 
14'h3daf : LOC =         127'b0000000000000000001000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000; // D (0x00001000000000020000000000000000) 
14'h06bc : LOC =         127'b0000000000000000010000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000; // D (0x00002000000000020000000000000000) 
14'h33ed : LOC =         127'b0000000000000000100000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000; // D (0x00004000000000020000000000000000) 
14'h1a38 : LOC =         127'b0000000000000001000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000; // D (0x00008000000000020000000000000000) 
14'h0ae5 : LOC =         127'b0000000000000010000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000; // D (0x00010000000000020000000000000000) 
14'h2b5f : LOC =         127'b0000000000000100000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000; // D (0x00020000000000020000000000000000) 
14'h2b5c : LOC =         127'b0000000000001000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000; // D (0x00040000000000020000000000000000) 
14'h2b5a : LOC =         127'b0000000000010000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000; // D (0x00080000000000020000000000000000) 
14'h2b56 : LOC =         127'b0000000000100000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000; // D (0x00100000000000020000000000000000) 
14'h2b4e : LOC =         127'b0000000001000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000; // D (0x00200000000000020000000000000000) 
14'h2b7e : LOC =         127'b0000000010000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000; // D (0x00400000000000020000000000000000) 
14'h2b1e : LOC =         127'b0000000100000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000; // D (0x00800000000000020000000000000000) 
14'h2bde : LOC =         127'b0000001000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000; // D (0x01000000000000020000000000000000) 
14'h2a5e : LOC =         127'b0000010000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000; // D (0x02000000000000020000000000000000) 
14'h295e : LOC =         127'b0000100000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000; // D (0x04000000000000020000000000000000) 
14'h2f5e : LOC =         127'b0001000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000; // D (0x08000000000000020000000000000000) 
14'h235e : LOC =         127'b0010000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000; // D (0x10000000000000020000000000000000) 
14'h3b5e : LOC =         127'b0100000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000; // D (0x20000000000000020000000000000000) 
14'h0b5e : LOC =         127'b1000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000; // D (0x40000000000000020000000000000000) 
14'h15cb : LOC =         127'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000; // S (0x00000000000000040000000000000000) 
14'h3e5d : LOC =         127'b0000000000000000000000000000000000000000000000000000000000011000000000000000000000000000000000000000000000000000000000000000000; // D (0x000000000000000c0000000000000000) 
14'h0190 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000101000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000000140000000000000000) 
14'h3d7d : LOC =         127'b0000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000000240000000000000000) 
14'h07d0 : LOC =         127'b0000000000000000000000000000000000000000000000000000000010001000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000000440000000000000000) 
14'h31fd : LOC =         127'b0000000000000000000000000000000000000000000000000000000100001000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000000840000000000000000) 
14'h1ed0 : LOC =         127'b0000000000000000000000000000000000000000000000000000001000001000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000001040000000000000000) 
14'h03fd : LOC =         127'b0000000000000000000000000000000000000000000000000000010000001000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000002040000000000000000) 
14'h39a7 : LOC =         127'b0000000000000000000000000000000000000000000000000000100000001000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000004040000000000000000) 
14'h0e64 : LOC =         127'b0000000000000000000000000000000000000000000000000001000000001000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000008040000000000000000) 
14'h2295 : LOC =         127'b0000000000000000000000000000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000010040000000000000000) 
14'h3800 : LOC =         127'b0000000000000000000000000000000000000000000000000100000000001000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000020040000000000000000) 
14'h0d2a : LOC =         127'b0000000000000000000000000000000000000000000000001000000000001000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000040040000000000000000) 
14'h2409 : LOC =         127'b0000000000000000000000000000000000000000000000010000000000001000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000080040000000000000000) 
14'h3538 : LOC =         127'b0000000000000000000000000000000000000000000000100000000000001000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000100040000000000000000) 
14'h175a : LOC =         127'b0000000000000000000000000000000000000000000001000000000000001000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000200040000000000000000) 
14'h10e9 : LOC =         127'b0000000000000000000000000000000000000000000010000000000000001000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000400040000000000000000) 
14'h1f8f : LOC =         127'b0000000000000000000000000000000000000000000100000000000000001000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000800040000000000000000) 
14'h0143 : LOC =         127'b0000000000000000000000000000000000000000001000000000000000001000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000001000040000000000000000) 
14'h3cdb : LOC =         127'b0000000000000000000000000000000000000000010000000000000000001000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000002000040000000000000000) 
14'h049c : LOC =         127'b0000000000000000000000000000000000000000100000000000000000001000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000004000040000000000000000) 
14'h3765 : LOC =         127'b0000000000000000000000000000000000000001000000000000000000001000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000008000040000000000000000) 
14'h13e0 : LOC =         127'b0000000000000000000000000000000000000010000000000000000000001000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000010000040000000000000000) 
14'h199d : LOC =         127'b0000000000000000000000000000000000000100000000000000000000001000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000020000040000000000000000) 
14'h0d67 : LOC =         127'b0000000000000000000000000000000000001000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000040000040000000000000000) 
14'h2493 : LOC =         127'b0000000000000000000000000000000000010000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000080000040000000000000000) 
14'h340c : LOC =         127'b0000000000000000000000000000000000100000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000100000040000000000000000) 
14'h1532 : LOC =         127'b0000000000000000000000000000000001000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000200000040000000000000000) 
14'h1439 : LOC =         127'b0000000000000000000000000000000010000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000400000040000000000000000) 
14'h162f : LOC =         127'b0000000000000000000000000000000100000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000800000040000000000000000) 
14'h1203 : LOC =         127'b0000000000000000000000000000001000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000001000000040000000000000000) 
14'h1a5b : LOC =         127'b0000000000000000000000000000010000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000002000000040000000000000000) 
14'h0aeb : LOC =         127'b0000000000000000000000000000100000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000004000000040000000000000000) 
14'h2b8b : LOC =         127'b0000000000000000000000000001000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000008000000040000000000000000) 
14'h2a3c : LOC =         127'b0000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000010000000040000000000000000) 
14'h2952 : LOC =         127'b0000000000000000000000000100000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000020000000040000000000000000) 
14'h2f8e : LOC =         127'b0000000000000000000000001000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000040000000040000000000000000) 
14'h2236 : LOC =         127'b0000000000000000000000010000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000080000000040000000000000000) 
14'h3946 : LOC =         127'b0000000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000100000000040000000000000000) 
14'h0fa6 : LOC =         127'b0000000000000000000001000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000200000000040000000000000000) 
14'h2111 : LOC =         127'b0000000000000000000010000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000400000000040000000000000000) 
14'h3f08 : LOC =         127'b0000000000000000000100000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000800000000040000000000000000) 
14'h033a : LOC =         127'b0000000000000000001000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000; // D (0x00001000000000040000000000000000) 
14'h3829 : LOC =         127'b0000000000000000010000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000; // D (0x00002000000000040000000000000000) 
14'h0d78 : LOC =         127'b0000000000000000100000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000; // D (0x00004000000000040000000000000000) 
14'h24ad : LOC =         127'b0000000000000001000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000; // D (0x00008000000000040000000000000000) 
14'h3470 : LOC =         127'b0000000000000010000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000; // D (0x00010000000000040000000000000000) 
14'h15ca : LOC =         127'b0000000000000100000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000; // D (0x00020000000000040000000000000000) 
14'h15c9 : LOC =         127'b0000000000001000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000; // D (0x00040000000000040000000000000000) 
14'h15cf : LOC =         127'b0000000000010000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000; // D (0x00080000000000040000000000000000) 
14'h15c3 : LOC =         127'b0000000000100000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000; // D (0x00100000000000040000000000000000) 
14'h15db : LOC =         127'b0000000001000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000; // D (0x00200000000000040000000000000000) 
14'h15eb : LOC =         127'b0000000010000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000; // D (0x00400000000000040000000000000000) 
14'h158b : LOC =         127'b0000000100000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000; // D (0x00800000000000040000000000000000) 
14'h154b : LOC =         127'b0000001000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000; // D (0x01000000000000040000000000000000) 
14'h14cb : LOC =         127'b0000010000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000; // D (0x02000000000000040000000000000000) 
14'h17cb : LOC =         127'b0000100000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000; // D (0x04000000000000040000000000000000) 
14'h11cb : LOC =         127'b0001000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000; // D (0x08000000000000040000000000000000) 
14'h1dcb : LOC =         127'b0010000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000; // D (0x10000000000000040000000000000000) 
14'h05cb : LOC =         127'b0100000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000; // D (0x20000000000000040000000000000000) 
14'h35cb : LOC =         127'b1000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000; // D (0x40000000000000040000000000000000) 
14'h2b96 : LOC =         127'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000; // S (0x00000000000000080000000000000000) 
14'h3fcd : LOC =         127'b0000000000000000000000000000000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000000180000000000000000) 
14'h0320 : LOC =         127'b0000000000000000000000000000000000000000000000000000000001010000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000000280000000000000000) 
14'h398d : LOC =         127'b0000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000000480000000000000000) 
14'h0fa0 : LOC =         127'b0000000000000000000000000000000000000000000000000000000100010000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000000880000000000000000) 
14'h208d : LOC =         127'b0000000000000000000000000000000000000000000000000000001000010000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000001080000000000000000) 
14'h3da0 : LOC =         127'b0000000000000000000000000000000000000000000000000000010000010000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000002080000000000000000) 
14'h07fa : LOC =         127'b0000000000000000000000000000000000000000000000000000100000010000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000004080000000000000000) 
14'h3039 : LOC =         127'b0000000000000000000000000000000000000000000000000001000000010000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000008080000000000000000) 
14'h1cc8 : LOC =         127'b0000000000000000000000000000000000000000000000000010000000010000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000010080000000000000000) 
14'h065d : LOC =         127'b0000000000000000000000000000000000000000000000000100000000010000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000020080000000000000000) 
14'h3377 : LOC =         127'b0000000000000000000000000000000000000000000000001000000000010000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000040080000000000000000) 
14'h1a54 : LOC =         127'b0000000000000000000000000000000000000000000000010000000000010000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000080080000000000000000) 
14'h0b65 : LOC =         127'b0000000000000000000000000000000000000000000000100000000000010000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000100080000000000000000) 
14'h2907 : LOC =         127'b0000000000000000000000000000000000000000000001000000000000010000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000200080000000000000000) 
14'h2eb4 : LOC =         127'b0000000000000000000000000000000000000000000010000000000000010000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000400080000000000000000) 
14'h21d2 : LOC =         127'b0000000000000000000000000000000000000000000100000000000000010000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000800080000000000000000) 
14'h3f1e : LOC =         127'b0000000000000000000000000000000000000000001000000000000000010000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000001000080000000000000000) 
14'h0286 : LOC =         127'b0000000000000000000000000000000000000000010000000000000000010000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000002000080000000000000000) 
14'h3ac1 : LOC =         127'b0000000000000000000000000000000000000000100000000000000000010000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000004000080000000000000000) 
14'h0938 : LOC =         127'b0000000000000000000000000000000000000001000000000000000000010000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000008000080000000000000000) 
14'h2dbd : LOC =         127'b0000000000000000000000000000000000000010000000000000000000010000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000010000080000000000000000) 
14'h27c0 : LOC =         127'b0000000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000020000080000000000000000) 
14'h333a : LOC =         127'b0000000000000000000000000000000000001000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000040000080000000000000000) 
14'h1ace : LOC =         127'b0000000000000000000000000000000000010000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000080000080000000000000000) 
14'h0a51 : LOC =         127'b0000000000000000000000000000000000100000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000100000080000000000000000) 
14'h2b6f : LOC =         127'b0000000000000000000000000000000001000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000200000080000000000000000) 
14'h2a64 : LOC =         127'b0000000000000000000000000000000010000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000400000080000000000000000) 
14'h2872 : LOC =         127'b0000000000000000000000000000000100000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000800000080000000000000000) 
14'h2c5e : LOC =         127'b0000000000000000000000000000001000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000001000000080000000000000000) 
14'h2406 : LOC =         127'b0000000000000000000000000000010000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000002000000080000000000000000) 
14'h34b6 : LOC =         127'b0000000000000000000000000000100000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000004000000080000000000000000) 
14'h15d6 : LOC =         127'b0000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000008000000080000000000000000) 
14'h1461 : LOC =         127'b0000000000000000000000000010000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000010000000080000000000000000) 
14'h170f : LOC =         127'b0000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000020000000080000000000000000) 
14'h11d3 : LOC =         127'b0000000000000000000000001000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000040000000080000000000000000) 
14'h1c6b : LOC =         127'b0000000000000000000000010000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000080000000080000000000000000) 
14'h071b : LOC =         127'b0000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000100000000080000000000000000) 
14'h31fb : LOC =         127'b0000000000000000000001000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000200000000080000000000000000) 
14'h1f4c : LOC =         127'b0000000000000000000010000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000400000000080000000000000000) 
14'h0155 : LOC =         127'b0000000000000000000100000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000800000000080000000000000000) 
14'h3d67 : LOC =         127'b0000000000000000001000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000; // D (0x00001000000000080000000000000000) 
14'h0674 : LOC =         127'b0000000000000000010000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000; // D (0x00002000000000080000000000000000) 
14'h3325 : LOC =         127'b0000000000000000100000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000; // D (0x00004000000000080000000000000000) 
14'h1af0 : LOC =         127'b0000000000000001000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000; // D (0x00008000000000080000000000000000) 
14'h0a2d : LOC =         127'b0000000000000010000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000; // D (0x00010000000000080000000000000000) 
14'h2b97 : LOC =         127'b0000000000000100000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000; // D (0x00020000000000080000000000000000) 
14'h2b94 : LOC =         127'b0000000000001000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000; // D (0x00040000000000080000000000000000) 
14'h2b92 : LOC =         127'b0000000000010000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000; // D (0x00080000000000080000000000000000) 
14'h2b9e : LOC =         127'b0000000000100000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000; // D (0x00100000000000080000000000000000) 
14'h2b86 : LOC =         127'b0000000001000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000; // D (0x00200000000000080000000000000000) 
14'h2bb6 : LOC =         127'b0000000010000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000; // D (0x00400000000000080000000000000000) 
14'h2bd6 : LOC =         127'b0000000100000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000; // D (0x00800000000000080000000000000000) 
14'h2b16 : LOC =         127'b0000001000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000; // D (0x01000000000000080000000000000000) 
14'h2a96 : LOC =         127'b0000010000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000; // D (0x02000000000000080000000000000000) 
14'h2996 : LOC =         127'b0000100000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000; // D (0x04000000000000080000000000000000) 
14'h2f96 : LOC =         127'b0001000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000; // D (0x08000000000000080000000000000000) 
14'h2396 : LOC =         127'b0010000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000; // D (0x10000000000000080000000000000000) 
14'h3b96 : LOC =         127'b0100000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000; // D (0x20000000000000080000000000000000) 
14'h0b96 : LOC =         127'b1000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000; // D (0x40000000000000080000000000000000) 
14'h145b : LOC =         127'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000; // S (0x00000000000000100000000000000000) 
14'h3ced : LOC =         127'b0000000000000000000000000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000000300000000000000000) 
14'h0640 : LOC =         127'b0000000000000000000000000000000000000000000000000000000010100000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000000500000000000000000) 
14'h306d : LOC =         127'b0000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000000900000000000000000) 
14'h1f40 : LOC =         127'b0000000000000000000000000000000000000000000000000000001000100000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000001100000000000000000) 
14'h026d : LOC =         127'b0000000000000000000000000000000000000000000000000000010000100000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000002100000000000000000) 
14'h3837 : LOC =         127'b0000000000000000000000000000000000000000000000000000100000100000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000004100000000000000000) 
14'h0ff4 : LOC =         127'b0000000000000000000000000000000000000000000000000001000000100000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000008100000000000000000) 
14'h2305 : LOC =         127'b0000000000000000000000000000000000000000000000000010000000100000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000010100000000000000000) 
14'h3990 : LOC =         127'b0000000000000000000000000000000000000000000000000100000000100000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000020100000000000000000) 
14'h0cba : LOC =         127'b0000000000000000000000000000000000000000000000001000000000100000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000040100000000000000000) 
14'h2599 : LOC =         127'b0000000000000000000000000000000000000000000000010000000000100000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000080100000000000000000) 
14'h34a8 : LOC =         127'b0000000000000000000000000000000000000000000000100000000000100000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000100100000000000000000) 
14'h16ca : LOC =         127'b0000000000000000000000000000000000000000000001000000000000100000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000200100000000000000000) 
14'h1179 : LOC =         127'b0000000000000000000000000000000000000000000010000000000000100000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000400100000000000000000) 
14'h1e1f : LOC =         127'b0000000000000000000000000000000000000000000100000000000000100000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000800100000000000000000) 
14'h00d3 : LOC =         127'b0000000000000000000000000000000000000000001000000000000000100000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000001000100000000000000000) 
14'h3d4b : LOC =         127'b0000000000000000000000000000000000000000010000000000000000100000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000002000100000000000000000) 
14'h050c : LOC =         127'b0000000000000000000000000000000000000000100000000000000000100000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000004000100000000000000000) 
14'h36f5 : LOC =         127'b0000000000000000000000000000000000000001000000000000000000100000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000008000100000000000000000) 
14'h1270 : LOC =         127'b0000000000000000000000000000000000000010000000000000000000100000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000010000100000000000000000) 
14'h180d : LOC =         127'b0000000000000000000000000000000000000100000000000000000000100000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000020000100000000000000000) 
14'h0cf7 : LOC =         127'b0000000000000000000000000000000000001000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000040000100000000000000000) 
14'h2503 : LOC =         127'b0000000000000000000000000000000000010000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000080000100000000000000000) 
14'h359c : LOC =         127'b0000000000000000000000000000000000100000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000100000100000000000000000) 
14'h14a2 : LOC =         127'b0000000000000000000000000000000001000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000200000100000000000000000) 
14'h15a9 : LOC =         127'b0000000000000000000000000000000010000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000400000100000000000000000) 
14'h17bf : LOC =         127'b0000000000000000000000000000000100000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000800000100000000000000000) 
14'h1393 : LOC =         127'b0000000000000000000000000000001000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000001000000100000000000000000) 
14'h1bcb : LOC =         127'b0000000000000000000000000000010000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000002000000100000000000000000) 
14'h0b7b : LOC =         127'b0000000000000000000000000000100000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000004000000100000000000000000) 
14'h2a1b : LOC =         127'b0000000000000000000000000001000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000008000000100000000000000000) 
14'h2bac : LOC =         127'b0000000000000000000000000010000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000010000000100000000000000000) 
14'h28c2 : LOC =         127'b0000000000000000000000000100000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000020000000100000000000000000) 
14'h2e1e : LOC =         127'b0000000000000000000000001000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000040000000100000000000000000) 
14'h23a6 : LOC =         127'b0000000000000000000000010000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000080000000100000000000000000) 
14'h38d6 : LOC =         127'b0000000000000000000000100000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000100000000100000000000000000) 
14'h0e36 : LOC =         127'b0000000000000000000001000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000200000000100000000000000000) 
14'h2081 : LOC =         127'b0000000000000000000010000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000400000000100000000000000000) 
14'h3e98 : LOC =         127'b0000000000000000000100000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000800000000100000000000000000) 
14'h02aa : LOC =         127'b0000000000000000001000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000; // D (0x00001000000000100000000000000000) 
14'h39b9 : LOC =         127'b0000000000000000010000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000; // D (0x00002000000000100000000000000000) 
14'h0ce8 : LOC =         127'b0000000000000000100000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000; // D (0x00004000000000100000000000000000) 
14'h253d : LOC =         127'b0000000000000001000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000; // D (0x00008000000000100000000000000000) 
14'h35e0 : LOC =         127'b0000000000000010000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000; // D (0x00010000000000100000000000000000) 
14'h145a : LOC =         127'b0000000000000100000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000; // D (0x00020000000000100000000000000000) 
14'h1459 : LOC =         127'b0000000000001000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000; // D (0x00040000000000100000000000000000) 
14'h145f : LOC =         127'b0000000000010000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000; // D (0x00080000000000100000000000000000) 
14'h1453 : LOC =         127'b0000000000100000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000; // D (0x00100000000000100000000000000000) 
14'h144b : LOC =         127'b0000000001000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000; // D (0x00200000000000100000000000000000) 
14'h147b : LOC =         127'b0000000010000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000; // D (0x00400000000000100000000000000000) 
14'h141b : LOC =         127'b0000000100000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000; // D (0x00800000000000100000000000000000) 
14'h14db : LOC =         127'b0000001000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000; // D (0x01000000000000100000000000000000) 
14'h155b : LOC =         127'b0000010000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000; // D (0x02000000000000100000000000000000) 
14'h165b : LOC =         127'b0000100000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000; // D (0x04000000000000100000000000000000) 
14'h105b : LOC =         127'b0001000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000; // D (0x08000000000000100000000000000000) 
14'h1c5b : LOC =         127'b0010000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000; // D (0x10000000000000100000000000000000) 
14'h045b : LOC =         127'b0100000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000; // D (0x20000000000000100000000000000000) 
14'h345b : LOC =         127'b1000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000; // D (0x40000000000000100000000000000000) 
14'h28b6 : LOC =         127'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000; // S (0x00000000000000200000000000000000) 
14'h3aad : LOC =         127'b0000000000000000000000000000000000000000000000000000000011000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000000600000000000000000) 
14'h0c80 : LOC =         127'b0000000000000000000000000000000000000000000000000000000101000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000000a00000000000000000) 
14'h23ad : LOC =         127'b0000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000001200000000000000000) 
14'h3e80 : LOC =         127'b0000000000000000000000000000000000000000000000000000010001000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000002200000000000000000) 
14'h04da : LOC =         127'b0000000000000000000000000000000000000000000000000000100001000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000004200000000000000000) 
14'h3319 : LOC =         127'b0000000000000000000000000000000000000000000000000001000001000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000008200000000000000000) 
14'h1fe8 : LOC =         127'b0000000000000000000000000000000000000000000000000010000001000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000010200000000000000000) 
14'h057d : LOC =         127'b0000000000000000000000000000000000000000000000000100000001000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000020200000000000000000) 
14'h3057 : LOC =         127'b0000000000000000000000000000000000000000000000001000000001000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000040200000000000000000) 
14'h1974 : LOC =         127'b0000000000000000000000000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000080200000000000000000) 
14'h0845 : LOC =         127'b0000000000000000000000000000000000000000000000100000000001000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000100200000000000000000) 
14'h2a27 : LOC =         127'b0000000000000000000000000000000000000000000001000000000001000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000200200000000000000000) 
14'h2d94 : LOC =         127'b0000000000000000000000000000000000000000000010000000000001000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000400200000000000000000) 
14'h22f2 : LOC =         127'b0000000000000000000000000000000000000000000100000000000001000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000800200000000000000000) 
14'h3c3e : LOC =         127'b0000000000000000000000000000000000000000001000000000000001000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000001000200000000000000000) 
14'h01a6 : LOC =         127'b0000000000000000000000000000000000000000010000000000000001000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000002000200000000000000000) 
14'h39e1 : LOC =         127'b0000000000000000000000000000000000000000100000000000000001000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000004000200000000000000000) 
14'h0a18 : LOC =         127'b0000000000000000000000000000000000000001000000000000000001000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000008000200000000000000000) 
14'h2e9d : LOC =         127'b0000000000000000000000000000000000000010000000000000000001000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000010000200000000000000000) 
14'h24e0 : LOC =         127'b0000000000000000000000000000000000000100000000000000000001000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000020000200000000000000000) 
14'h301a : LOC =         127'b0000000000000000000000000000000000001000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000040000200000000000000000) 
14'h19ee : LOC =         127'b0000000000000000000000000000000000010000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000080000200000000000000000) 
14'h0971 : LOC =         127'b0000000000000000000000000000000000100000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000100000200000000000000000) 
14'h284f : LOC =         127'b0000000000000000000000000000000001000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000200000200000000000000000) 
14'h2944 : LOC =         127'b0000000000000000000000000000000010000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000400000200000000000000000) 
14'h2b52 : LOC =         127'b0000000000000000000000000000000100000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000800000200000000000000000) 
14'h2f7e : LOC =         127'b0000000000000000000000000000001000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000001000000200000000000000000) 
14'h2726 : LOC =         127'b0000000000000000000000000000010000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000002000000200000000000000000) 
14'h3796 : LOC =         127'b0000000000000000000000000000100000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000004000000200000000000000000) 
14'h16f6 : LOC =         127'b0000000000000000000000000001000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000008000000200000000000000000) 
14'h1741 : LOC =         127'b0000000000000000000000000010000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000010000000200000000000000000) 
14'h142f : LOC =         127'b0000000000000000000000000100000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000020000000200000000000000000) 
14'h12f3 : LOC =         127'b0000000000000000000000001000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000040000000200000000000000000) 
14'h1f4b : LOC =         127'b0000000000000000000000010000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000080000000200000000000000000) 
14'h043b : LOC =         127'b0000000000000000000000100000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000100000000200000000000000000) 
14'h32db : LOC =         127'b0000000000000000000001000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000200000000200000000000000000) 
14'h1c6c : LOC =         127'b0000000000000000000010000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000400000000200000000000000000) 
14'h0275 : LOC =         127'b0000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000800000000200000000000000000) 
14'h3e47 : LOC =         127'b0000000000000000001000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00001000000000200000000000000000) 
14'h0554 : LOC =         127'b0000000000000000010000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00002000000000200000000000000000) 
14'h3005 : LOC =         127'b0000000000000000100000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00004000000000200000000000000000) 
14'h19d0 : LOC =         127'b0000000000000001000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00008000000000200000000000000000) 
14'h090d : LOC =         127'b0000000000000010000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00010000000000200000000000000000) 
14'h28b7 : LOC =         127'b0000000000000100000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00020000000000200000000000000000) 
14'h28b4 : LOC =         127'b0000000000001000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00040000000000200000000000000000) 
14'h28b2 : LOC =         127'b0000000000010000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00080000000000200000000000000000) 
14'h28be : LOC =         127'b0000000000100000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00100000000000200000000000000000) 
14'h28a6 : LOC =         127'b0000000001000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00200000000000200000000000000000) 
14'h2896 : LOC =         127'b0000000010000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00400000000000200000000000000000) 
14'h28f6 : LOC =         127'b0000000100000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00800000000000200000000000000000) 
14'h2836 : LOC =         127'b0000001000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000; // D (0x01000000000000200000000000000000) 
14'h29b6 : LOC =         127'b0000010000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000; // D (0x02000000000000200000000000000000) 
14'h2ab6 : LOC =         127'b0000100000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000; // D (0x04000000000000200000000000000000) 
14'h2cb6 : LOC =         127'b0001000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000; // D (0x08000000000000200000000000000000) 
14'h20b6 : LOC =         127'b0010000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000; // D (0x10000000000000200000000000000000) 
14'h38b6 : LOC =         127'b0100000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000; // D (0x20000000000000200000000000000000) 
14'h08b6 : LOC =         127'b1000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000; // D (0x40000000000000200000000000000000) 
14'h121b : LOC =         127'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000; // S (0x00000000000000400000000000000000) 
14'h362d : LOC =         127'b0000000000000000000000000000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000000c00000000000000000) 
14'h1900 : LOC =         127'b0000000000000000000000000000000000000000000000000000001010000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000001400000000000000000) 
14'h042d : LOC =         127'b0000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000002400000000000000000) 
14'h3e77 : LOC =         127'b0000000000000000000000000000000000000000000000000000100010000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000004400000000000000000) 
14'h09b4 : LOC =         127'b0000000000000000000000000000000000000000000000000001000010000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000008400000000000000000) 
14'h2545 : LOC =         127'b0000000000000000000000000000000000000000000000000010000010000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000010400000000000000000) 
14'h3fd0 : LOC =         127'b0000000000000000000000000000000000000000000000000100000010000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000020400000000000000000) 
14'h0afa : LOC =         127'b0000000000000000000000000000000000000000000000001000000010000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000040400000000000000000) 
14'h23d9 : LOC =         127'b0000000000000000000000000000000000000000000000010000000010000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000080400000000000000000) 
14'h32e8 : LOC =         127'b0000000000000000000000000000000000000000000000100000000010000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000100400000000000000000) 
14'h108a : LOC =         127'b0000000000000000000000000000000000000000000001000000000010000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000200400000000000000000) 
14'h1739 : LOC =         127'b0000000000000000000000000000000000000000000010000000000010000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000400400000000000000000) 
14'h185f : LOC =         127'b0000000000000000000000000000000000000000000100000000000010000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000800400000000000000000) 
14'h0693 : LOC =         127'b0000000000000000000000000000000000000000001000000000000010000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000001000400000000000000000) 
14'h3b0b : LOC =         127'b0000000000000000000000000000000000000000010000000000000010000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000002000400000000000000000) 
14'h034c : LOC =         127'b0000000000000000000000000000000000000000100000000000000010000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000004000400000000000000000) 
14'h30b5 : LOC =         127'b0000000000000000000000000000000000000001000000000000000010000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000008000400000000000000000) 
14'h1430 : LOC =         127'b0000000000000000000000000000000000000010000000000000000010000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000010000400000000000000000) 
14'h1e4d : LOC =         127'b0000000000000000000000000000000000000100000000000000000010000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000020000400000000000000000) 
14'h0ab7 : LOC =         127'b0000000000000000000000000000000000001000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000040000400000000000000000) 
14'h2343 : LOC =         127'b0000000000000000000000000000000000010000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000080000400000000000000000) 
14'h33dc : LOC =         127'b0000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000100000400000000000000000) 
14'h12e2 : LOC =         127'b0000000000000000000000000000000001000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000200000400000000000000000) 
14'h13e9 : LOC =         127'b0000000000000000000000000000000010000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000400000400000000000000000) 
14'h11ff : LOC =         127'b0000000000000000000000000000000100000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000800000400000000000000000) 
14'h15d3 : LOC =         127'b0000000000000000000000000000001000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000001000000400000000000000000) 
14'h1d8b : LOC =         127'b0000000000000000000000000000010000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000002000000400000000000000000) 
14'h0d3b : LOC =         127'b0000000000000000000000000000100000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000004000000400000000000000000) 
14'h2c5b : LOC =         127'b0000000000000000000000000001000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000008000000400000000000000000) 
14'h2dec : LOC =         127'b0000000000000000000000000010000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000010000000400000000000000000) 
14'h2e82 : LOC =         127'b0000000000000000000000000100000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000020000000400000000000000000) 
14'h285e : LOC =         127'b0000000000000000000000001000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000040000000400000000000000000) 
14'h25e6 : LOC =         127'b0000000000000000000000010000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000080000000400000000000000000) 
14'h3e96 : LOC =         127'b0000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000100000000400000000000000000) 
14'h0876 : LOC =         127'b0000000000000000000001000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000200000000400000000000000000) 
14'h26c1 : LOC =         127'b0000000000000000000010000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000400000000400000000000000000) 
14'h38d8 : LOC =         127'b0000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000800000000400000000000000000) 
14'h04ea : LOC =         127'b0000000000000000001000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00001000000000400000000000000000) 
14'h3ff9 : LOC =         127'b0000000000000000010000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00002000000000400000000000000000) 
14'h0aa8 : LOC =         127'b0000000000000000100000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00004000000000400000000000000000) 
14'h237d : LOC =         127'b0000000000000001000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00008000000000400000000000000000) 
14'h33a0 : LOC =         127'b0000000000000010000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00010000000000400000000000000000) 
14'h121a : LOC =         127'b0000000000000100000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00020000000000400000000000000000) 
14'h1219 : LOC =         127'b0000000000001000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00040000000000400000000000000000) 
14'h121f : LOC =         127'b0000000000010000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00080000000000400000000000000000) 
14'h1213 : LOC =         127'b0000000000100000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00100000000000400000000000000000) 
14'h120b : LOC =         127'b0000000001000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00200000000000400000000000000000) 
14'h123b : LOC =         127'b0000000010000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00400000000000400000000000000000) 
14'h125b : LOC =         127'b0000000100000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00800000000000400000000000000000) 
14'h129b : LOC =         127'b0000001000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000; // D (0x01000000000000400000000000000000) 
14'h131b : LOC =         127'b0000010000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000; // D (0x02000000000000400000000000000000) 
14'h101b : LOC =         127'b0000100000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000; // D (0x04000000000000400000000000000000) 
14'h161b : LOC =         127'b0001000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000; // D (0x08000000000000400000000000000000) 
14'h1a1b : LOC =         127'b0010000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000; // D (0x10000000000000400000000000000000) 
14'h021b : LOC =         127'b0100000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000; // D (0x20000000000000400000000000000000) 
14'h321b : LOC =         127'b1000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000; // D (0x40000000000000400000000000000000) 
14'h2436 : LOC =         127'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000; // S (0x00000000000000800000000000000000) 
14'h2f2d : LOC =         127'b0000000000000000000000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000001800000000000000000) 
14'h3200 : LOC =         127'b0000000000000000000000000000000000000000000000000000010100000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000002800000000000000000) 
14'h085a : LOC =         127'b0000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000004800000000000000000) 
14'h3f99 : LOC =         127'b0000000000000000000000000000000000000000000000000001000100000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000008800000000000000000) 
14'h1368 : LOC =         127'b0000000000000000000000000000000000000000000000000010000100000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000010800000000000000000) 
14'h09fd : LOC =         127'b0000000000000000000000000000000000000000000000000100000100000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000020800000000000000000) 
14'h3cd7 : LOC =         127'b0000000000000000000000000000000000000000000000001000000100000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000040800000000000000000) 
14'h15f4 : LOC =         127'b0000000000000000000000000000000000000000000000010000000100000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000080800000000000000000) 
14'h04c5 : LOC =         127'b0000000000000000000000000000000000000000000000100000000100000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000100800000000000000000) 
14'h26a7 : LOC =         127'b0000000000000000000000000000000000000000000001000000000100000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000200800000000000000000) 
14'h2114 : LOC =         127'b0000000000000000000000000000000000000000000010000000000100000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000400800000000000000000) 
14'h2e72 : LOC =         127'b0000000000000000000000000000000000000000000100000000000100000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000800800000000000000000) 
14'h30be : LOC =         127'b0000000000000000000000000000000000000000001000000000000100000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000001000800000000000000000) 
14'h0d26 : LOC =         127'b0000000000000000000000000000000000000000010000000000000100000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000002000800000000000000000) 
14'h3561 : LOC =         127'b0000000000000000000000000000000000000000100000000000000100000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000004000800000000000000000) 
14'h0698 : LOC =         127'b0000000000000000000000000000000000000001000000000000000100000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000008000800000000000000000) 
14'h221d : LOC =         127'b0000000000000000000000000000000000000010000000000000000100000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000010000800000000000000000) 
14'h2860 : LOC =         127'b0000000000000000000000000000000000000100000000000000000100000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000020000800000000000000000) 
14'h3c9a : LOC =         127'b0000000000000000000000000000000000001000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000040000800000000000000000) 
14'h156e : LOC =         127'b0000000000000000000000000000000000010000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000080000800000000000000000) 
14'h05f1 : LOC =         127'b0000000000000000000000000000000000100000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000100000800000000000000000) 
14'h24cf : LOC =         127'b0000000000000000000000000000000001000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000200000800000000000000000) 
14'h25c4 : LOC =         127'b0000000000000000000000000000000010000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000400000800000000000000000) 
14'h27d2 : LOC =         127'b0000000000000000000000000000000100000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000800000800000000000000000) 
14'h23fe : LOC =         127'b0000000000000000000000000000001000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000001000000800000000000000000) 
14'h2ba6 : LOC =         127'b0000000000000000000000000000010000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000002000000800000000000000000) 
14'h3b16 : LOC =         127'b0000000000000000000000000000100000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000004000000800000000000000000) 
14'h1a76 : LOC =         127'b0000000000000000000000000001000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000008000000800000000000000000) 
14'h1bc1 : LOC =         127'b0000000000000000000000000010000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000010000000800000000000000000) 
14'h18af : LOC =         127'b0000000000000000000000000100000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000020000000800000000000000000) 
14'h1e73 : LOC =         127'b0000000000000000000000001000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000040000000800000000000000000) 
14'h13cb : LOC =         127'b0000000000000000000000010000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000080000000800000000000000000) 
14'h08bb : LOC =         127'b0000000000000000000000100000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000100000000800000000000000000) 
14'h3e5b : LOC =         127'b0000000000000000000001000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000200000000800000000000000000) 
14'h10ec : LOC =         127'b0000000000000000000010000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000400000000800000000000000000) 
14'h0ef5 : LOC =         127'b0000000000000000000100000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000800000000800000000000000000) 
14'h32c7 : LOC =         127'b0000000000000000001000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00001000000000800000000000000000) 
14'h09d4 : LOC =         127'b0000000000000000010000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00002000000000800000000000000000) 
14'h3c85 : LOC =         127'b0000000000000000100000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00004000000000800000000000000000) 
14'h1550 : LOC =         127'b0000000000000001000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00008000000000800000000000000000) 
14'h058d : LOC =         127'b0000000000000010000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00010000000000800000000000000000) 
14'h2437 : LOC =         127'b0000000000000100000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00020000000000800000000000000000) 
14'h2434 : LOC =         127'b0000000000001000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00040000000000800000000000000000) 
14'h2432 : LOC =         127'b0000000000010000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00080000000000800000000000000000) 
14'h243e : LOC =         127'b0000000000100000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00100000000000800000000000000000) 
14'h2426 : LOC =         127'b0000000001000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00200000000000800000000000000000) 
14'h2416 : LOC =         127'b0000000010000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00400000000000800000000000000000) 
14'h2476 : LOC =         127'b0000000100000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00800000000000800000000000000000) 
14'h24b6 : LOC =         127'b0000001000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000; // D (0x01000000000000800000000000000000) 
14'h2536 : LOC =         127'b0000010000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000; // D (0x02000000000000800000000000000000) 
14'h2636 : LOC =         127'b0000100000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000; // D (0x04000000000000800000000000000000) 
14'h2036 : LOC =         127'b0001000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000; // D (0x08000000000000800000000000000000) 
14'h2c36 : LOC =         127'b0010000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000; // D (0x10000000000000800000000000000000) 
14'h3436 : LOC =         127'b0100000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000; // D (0x20000000000000800000000000000000) 
14'h0436 : LOC =         127'b1000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000; // D (0x40000000000000800000000000000000) 
14'h0b1b : LOC =         127'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000; // S (0x00000000000001000000000000000000) 
14'h1d2d : LOC =         127'b0000000000000000000000000000000000000000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000003000000000000000000) 
14'h2777 : LOC =         127'b0000000000000000000000000000000000000000000000000000101000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000005000000000000000000) 
14'h10b4 : LOC =         127'b0000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000009000000000000000000) 
14'h3c45 : LOC =         127'b0000000000000000000000000000000000000000000000000010001000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000011000000000000000000) 
14'h26d0 : LOC =         127'b0000000000000000000000000000000000000000000000000100001000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000021000000000000000000) 
14'h13fa : LOC =         127'b0000000000000000000000000000000000000000000000001000001000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000041000000000000000000) 
14'h3ad9 : LOC =         127'b0000000000000000000000000000000000000000000000010000001000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000081000000000000000000) 
14'h2be8 : LOC =         127'b0000000000000000000000000000000000000000000000100000001000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000101000000000000000000) 
14'h098a : LOC =         127'b0000000000000000000000000000000000000000000001000000001000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000201000000000000000000) 
14'h0e39 : LOC =         127'b0000000000000000000000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000401000000000000000000) 
14'h015f : LOC =         127'b0000000000000000000000000000000000000000000100000000001000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000801000000000000000000) 
14'h1f93 : LOC =         127'b0000000000000000000000000000000000000000001000000000001000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000001001000000000000000000) 
14'h220b : LOC =         127'b0000000000000000000000000000000000000000010000000000001000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000002001000000000000000000) 
14'h1a4c : LOC =         127'b0000000000000000000000000000000000000000100000000000001000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000004001000000000000000000) 
14'h29b5 : LOC =         127'b0000000000000000000000000000000000000001000000000000001000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000008001000000000000000000) 
14'h0d30 : LOC =         127'b0000000000000000000000000000000000000010000000000000001000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000010001000000000000000000) 
14'h074d : LOC =         127'b0000000000000000000000000000000000000100000000000000001000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000020001000000000000000000) 
14'h13b7 : LOC =         127'b0000000000000000000000000000000000001000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000040001000000000000000000) 
14'h3a43 : LOC =         127'b0000000000000000000000000000000000010000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000080001000000000000000000) 
14'h2adc : LOC =         127'b0000000000000000000000000000000000100000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000100001000000000000000000) 
14'h0be2 : LOC =         127'b0000000000000000000000000000000001000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000200001000000000000000000) 
14'h0ae9 : LOC =         127'b0000000000000000000000000000000010000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000400001000000000000000000) 
14'h08ff : LOC =         127'b0000000000000000000000000000000100000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000800001000000000000000000) 
14'h0cd3 : LOC =         127'b0000000000000000000000000000001000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000001000001000000000000000000) 
14'h048b : LOC =         127'b0000000000000000000000000000010000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000002000001000000000000000000) 
14'h143b : LOC =         127'b0000000000000000000000000000100000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000004000001000000000000000000) 
14'h355b : LOC =         127'b0000000000000000000000000001000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000008000001000000000000000000) 
14'h34ec : LOC =         127'b0000000000000000000000000010000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000010000001000000000000000000) 
14'h3782 : LOC =         127'b0000000000000000000000000100000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000020000001000000000000000000) 
14'h315e : LOC =         127'b0000000000000000000000001000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000040000001000000000000000000) 
14'h3ce6 : LOC =         127'b0000000000000000000000010000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000080000001000000000000000000) 
14'h2796 : LOC =         127'b0000000000000000000000100000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000100000001000000000000000000) 
14'h1176 : LOC =         127'b0000000000000000000001000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000200000001000000000000000000) 
14'h3fc1 : LOC =         127'b0000000000000000000010000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000400000001000000000000000000) 
14'h21d8 : LOC =         127'b0000000000000000000100000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000800000001000000000000000000) 
14'h1dea : LOC =         127'b0000000000000000001000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00001000000001000000000000000000) 
14'h26f9 : LOC =         127'b0000000000000000010000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00002000000001000000000000000000) 
14'h13a8 : LOC =         127'b0000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00004000000001000000000000000000) 
14'h3a7d : LOC =         127'b0000000000000001000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00008000000001000000000000000000) 
14'h2aa0 : LOC =         127'b0000000000000010000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00010000000001000000000000000000) 
14'h0b1a : LOC =         127'b0000000000000100000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00020000000001000000000000000000) 
14'h0b19 : LOC =         127'b0000000000001000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00040000000001000000000000000000) 
14'h0b1f : LOC =         127'b0000000000010000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00080000000001000000000000000000) 
14'h0b13 : LOC =         127'b0000000000100000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00100000000001000000000000000000) 
14'h0b0b : LOC =         127'b0000000001000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00200000000001000000000000000000) 
14'h0b3b : LOC =         127'b0000000010000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00400000000001000000000000000000) 
14'h0b5b : LOC =         127'b0000000100000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00800000000001000000000000000000) 
14'h0b9b : LOC =         127'b0000001000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x01000000000001000000000000000000) 
14'h0a1b : LOC =         127'b0000010000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x02000000000001000000000000000000) 
14'h091b : LOC =         127'b0000100000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x04000000000001000000000000000000) 
14'h0f1b : LOC =         127'b0001000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x08000000000001000000000000000000) 
14'h031b : LOC =         127'b0010000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x10000000000001000000000000000000) 
14'h1b1b : LOC =         127'b0100000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x20000000000001000000000000000000) 
14'h2b1b : LOC =         127'b1000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x40000000000001000000000000000000) 
14'h1636 : LOC =         127'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000; // S (0x00000000000002000000000000000000) 
14'h3a5a : LOC =         127'b0000000000000000000000000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000006000000000000000000) 
14'h0d99 : LOC =         127'b0000000000000000000000000000000000000000000000000001010000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x0000000000000a000000000000000000) 
14'h2168 : LOC =         127'b0000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000012000000000000000000) 
14'h3bfd : LOC =         127'b0000000000000000000000000000000000000000000000000100010000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000022000000000000000000) 
14'h0ed7 : LOC =         127'b0000000000000000000000000000000000000000000000001000010000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000042000000000000000000) 
14'h27f4 : LOC =         127'b0000000000000000000000000000000000000000000000010000010000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000082000000000000000000) 
14'h36c5 : LOC =         127'b0000000000000000000000000000000000000000000000100000010000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000102000000000000000000) 
14'h14a7 : LOC =         127'b0000000000000000000000000000000000000000000001000000010000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000202000000000000000000) 
14'h1314 : LOC =         127'b0000000000000000000000000000000000000000000010000000010000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000402000000000000000000) 
14'h1c72 : LOC =         127'b0000000000000000000000000000000000000000000100000000010000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000802000000000000000000) 
14'h02be : LOC =         127'b0000000000000000000000000000000000000000001000000000010000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000001002000000000000000000) 
14'h3f26 : LOC =         127'b0000000000000000000000000000000000000000010000000000010000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000002002000000000000000000) 
14'h0761 : LOC =         127'b0000000000000000000000000000000000000000100000000000010000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000004002000000000000000000) 
14'h3498 : LOC =         127'b0000000000000000000000000000000000000001000000000000010000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000008002000000000000000000) 
14'h101d : LOC =         127'b0000000000000000000000000000000000000010000000000000010000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000010002000000000000000000) 
14'h1a60 : LOC =         127'b0000000000000000000000000000000000000100000000000000010000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000020002000000000000000000) 
14'h0e9a : LOC =         127'b0000000000000000000000000000000000001000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000040002000000000000000000) 
14'h276e : LOC =         127'b0000000000000000000000000000000000010000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000080002000000000000000000) 
14'h37f1 : LOC =         127'b0000000000000000000000000000000000100000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000100002000000000000000000) 
14'h16cf : LOC =         127'b0000000000000000000000000000000001000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000200002000000000000000000) 
14'h17c4 : LOC =         127'b0000000000000000000000000000000010000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000400002000000000000000000) 
14'h15d2 : LOC =         127'b0000000000000000000000000000000100000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000800002000000000000000000) 
14'h11fe : LOC =         127'b0000000000000000000000000000001000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000001000002000000000000000000) 
14'h19a6 : LOC =         127'b0000000000000000000000000000010000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000002000002000000000000000000) 
14'h0916 : LOC =         127'b0000000000000000000000000000100000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000004000002000000000000000000) 
14'h2876 : LOC =         127'b0000000000000000000000000001000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000008000002000000000000000000) 
14'h29c1 : LOC =         127'b0000000000000000000000000010000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000010000002000000000000000000) 
14'h2aaf : LOC =         127'b0000000000000000000000000100000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000020000002000000000000000000) 
14'h2c73 : LOC =         127'b0000000000000000000000001000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000040000002000000000000000000) 
14'h21cb : LOC =         127'b0000000000000000000000010000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000080000002000000000000000000) 
14'h3abb : LOC =         127'b0000000000000000000000100000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000100000002000000000000000000) 
14'h0c5b : LOC =         127'b0000000000000000000001000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000200000002000000000000000000) 
14'h22ec : LOC =         127'b0000000000000000000010000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000400000002000000000000000000) 
14'h3cf5 : LOC =         127'b0000000000000000000100000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000800000002000000000000000000) 
14'h00c7 : LOC =         127'b0000000000000000001000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00001000000002000000000000000000) 
14'h3bd4 : LOC =         127'b0000000000000000010000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00002000000002000000000000000000) 
14'h0e85 : LOC =         127'b0000000000000000100000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00004000000002000000000000000000) 
14'h2750 : LOC =         127'b0000000000000001000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00008000000002000000000000000000) 
14'h378d : LOC =         127'b0000000000000010000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00010000000002000000000000000000) 
14'h1637 : LOC =         127'b0000000000000100000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00020000000002000000000000000000) 
14'h1634 : LOC =         127'b0000000000001000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00040000000002000000000000000000) 
14'h1632 : LOC =         127'b0000000000010000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00080000000002000000000000000000) 
14'h163e : LOC =         127'b0000000000100000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00100000000002000000000000000000) 
14'h1626 : LOC =         127'b0000000001000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00200000000002000000000000000000) 
14'h1616 : LOC =         127'b0000000010000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00400000000002000000000000000000) 
14'h1676 : LOC =         127'b0000000100000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00800000000002000000000000000000) 
14'h16b6 : LOC =         127'b0000001000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x01000000000002000000000000000000) 
14'h1736 : LOC =         127'b0000010000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x02000000000002000000000000000000) 
14'h1436 : LOC =         127'b0000100000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x04000000000002000000000000000000) 
14'h1236 : LOC =         127'b0001000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x08000000000002000000000000000000) 
14'h1e36 : LOC =         127'b0010000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x10000000000002000000000000000000) 
14'h0636 : LOC =         127'b0100000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x20000000000002000000000000000000) 
14'h3636 : LOC =         127'b1000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x40000000000002000000000000000000) 
14'h2c6c : LOC =         127'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000; // S (0x00000000000004000000000000000000) 
14'h37c3 : LOC =         127'b0000000000000000000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x0000000000000c000000000000000000) 
14'h1b32 : LOC =         127'b0000000000000000000000000000000000000000000000000010100000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000014000000000000000000) 
14'h01a7 : LOC =         127'b0000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000024000000000000000000) 
14'h348d : LOC =         127'b0000000000000000000000000000000000000000000000001000100000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000044000000000000000000) 
14'h1dae : LOC =         127'b0000000000000000000000000000000000000000000000010000100000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000084000000000000000000) 
14'h0c9f : LOC =         127'b0000000000000000000000000000000000000000000000100000100000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000104000000000000000000) 
14'h2efd : LOC =         127'b0000000000000000000000000000000000000000000001000000100000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000204000000000000000000) 
14'h294e : LOC =         127'b0000000000000000000000000000000000000000000010000000100000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000404000000000000000000) 
14'h2628 : LOC =         127'b0000000000000000000000000000000000000000000100000000100000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000804000000000000000000) 
14'h38e4 : LOC =         127'b0000000000000000000000000000000000000000001000000000100000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000001004000000000000000000) 
14'h057c : LOC =         127'b0000000000000000000000000000000000000000010000000000100000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000002004000000000000000000) 
14'h3d3b : LOC =         127'b0000000000000000000000000000000000000000100000000000100000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000004004000000000000000000) 
14'h0ec2 : LOC =         127'b0000000000000000000000000000000000000001000000000000100000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000008004000000000000000000) 
14'h2a47 : LOC =         127'b0000000000000000000000000000000000000010000000000000100000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000010004000000000000000000) 
14'h203a : LOC =         127'b0000000000000000000000000000000000000100000000000000100000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000020004000000000000000000) 
14'h34c0 : LOC =         127'b0000000000000000000000000000000000001000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000040004000000000000000000) 
14'h1d34 : LOC =         127'b0000000000000000000000000000000000010000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000080004000000000000000000) 
14'h0dab : LOC =         127'b0000000000000000000000000000000000100000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000100004000000000000000000) 
14'h2c95 : LOC =         127'b0000000000000000000000000000000001000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000200004000000000000000000) 
14'h2d9e : LOC =         127'b0000000000000000000000000000000010000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000400004000000000000000000) 
14'h2f88 : LOC =         127'b0000000000000000000000000000000100000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000800004000000000000000000) 
14'h2ba4 : LOC =         127'b0000000000000000000000000000001000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000001000004000000000000000000) 
14'h23fc : LOC =         127'b0000000000000000000000000000010000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000002000004000000000000000000) 
14'h334c : LOC =         127'b0000000000000000000000000000100000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000004000004000000000000000000) 
14'h122c : LOC =         127'b0000000000000000000000000001000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000008000004000000000000000000) 
14'h139b : LOC =         127'b0000000000000000000000000010000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000010000004000000000000000000) 
14'h10f5 : LOC =         127'b0000000000000000000000000100000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000020000004000000000000000000) 
14'h1629 : LOC =         127'b0000000000000000000000001000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000040000004000000000000000000) 
14'h1b91 : LOC =         127'b0000000000000000000000010000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000080000004000000000000000000) 
14'h00e1 : LOC =         127'b0000000000000000000000100000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000100000004000000000000000000) 
14'h3601 : LOC =         127'b0000000000000000000001000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000200000004000000000000000000) 
14'h18b6 : LOC =         127'b0000000000000000000010000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000400000004000000000000000000) 
14'h06af : LOC =         127'b0000000000000000000100000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000800000004000000000000000000) 
14'h3a9d : LOC =         127'b0000000000000000001000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00001000000004000000000000000000) 
14'h018e : LOC =         127'b0000000000000000010000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00002000000004000000000000000000) 
14'h34df : LOC =         127'b0000000000000000100000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00004000000004000000000000000000) 
14'h1d0a : LOC =         127'b0000000000000001000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00008000000004000000000000000000) 
14'h0dd7 : LOC =         127'b0000000000000010000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00010000000004000000000000000000) 
14'h2c6d : LOC =         127'b0000000000000100000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00020000000004000000000000000000) 
14'h2c6e : LOC =         127'b0000000000001000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00040000000004000000000000000000) 
14'h2c68 : LOC =         127'b0000000000010000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00080000000004000000000000000000) 
14'h2c64 : LOC =         127'b0000000000100000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00100000000004000000000000000000) 
14'h2c7c : LOC =         127'b0000000001000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00200000000004000000000000000000) 
14'h2c4c : LOC =         127'b0000000010000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00400000000004000000000000000000) 
14'h2c2c : LOC =         127'b0000000100000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00800000000004000000000000000000) 
14'h2cec : LOC =         127'b0000001000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x01000000000004000000000000000000) 
14'h2d6c : LOC =         127'b0000010000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x02000000000004000000000000000000) 
14'h2e6c : LOC =         127'b0000100000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x04000000000004000000000000000000) 
14'h286c : LOC =         127'b0001000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x08000000000004000000000000000000) 
14'h246c : LOC =         127'b0010000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x10000000000004000000000000000000) 
14'h3c6c : LOC =         127'b0100000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x20000000000004000000000000000000) 
14'h0c6c : LOC =         127'b1000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x40000000000004000000000000000000) 
14'h1baf : LOC =         127'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000; // S (0x00000000000008000000000000000000) 
14'h2cf1 : LOC =         127'b0000000000000000000000000000000000000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000018000000000000000000) 
14'h3664 : LOC =         127'b0000000000000000000000000000000000000000000000000101000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000028000000000000000000) 
14'h034e : LOC =         127'b0000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000048000000000000000000) 
14'h2a6d : LOC =         127'b0000000000000000000000000000000000000000000000010001000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000088000000000000000000) 
14'h3b5c : LOC =         127'b0000000000000000000000000000000000000000000000100001000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000108000000000000000000) 
14'h193e : LOC =         127'b0000000000000000000000000000000000000000000001000001000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000208000000000000000000) 
14'h1e8d : LOC =         127'b0000000000000000000000000000000000000000000010000001000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000408000000000000000000) 
14'h11eb : LOC =         127'b0000000000000000000000000000000000000000000100000001000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000808000000000000000000) 
14'h0f27 : LOC =         127'b0000000000000000000000000000000000000000001000000001000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000001008000000000000000000) 
14'h32bf : LOC =         127'b0000000000000000000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000002008000000000000000000) 
14'h0af8 : LOC =         127'b0000000000000000000000000000000000000000100000000001000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000004008000000000000000000) 
14'h3901 : LOC =         127'b0000000000000000000000000000000000000001000000000001000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000008008000000000000000000) 
14'h1d84 : LOC =         127'b0000000000000000000000000000000000000010000000000001000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000010008000000000000000000) 
14'h17f9 : LOC =         127'b0000000000000000000000000000000000000100000000000001000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000020008000000000000000000) 
14'h0303 : LOC =         127'b0000000000000000000000000000000000001000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000040008000000000000000000) 
14'h2af7 : LOC =         127'b0000000000000000000000000000000000010000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000080008000000000000000000) 
14'h3a68 : LOC =         127'b0000000000000000000000000000000000100000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000100008000000000000000000) 
14'h1b56 : LOC =         127'b0000000000000000000000000000000001000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000200008000000000000000000) 
14'h1a5d : LOC =         127'b0000000000000000000000000000000010000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000400008000000000000000000) 
14'h184b : LOC =         127'b0000000000000000000000000000000100000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000800008000000000000000000) 
14'h1c67 : LOC =         127'b0000000000000000000000000000001000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000001000008000000000000000000) 
14'h143f : LOC =         127'b0000000000000000000000000000010000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000002000008000000000000000000) 
14'h048f : LOC =         127'b0000000000000000000000000000100000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000004000008000000000000000000) 
14'h25ef : LOC =         127'b0000000000000000000000000001000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000008000008000000000000000000) 
14'h2458 : LOC =         127'b0000000000000000000000000010000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000010000008000000000000000000) 
14'h2736 : LOC =         127'b0000000000000000000000000100000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000020000008000000000000000000) 
14'h21ea : LOC =         127'b0000000000000000000000001000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000040000008000000000000000000) 
14'h2c52 : LOC =         127'b0000000000000000000000010000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000080000008000000000000000000) 
14'h3722 : LOC =         127'b0000000000000000000000100000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000100000008000000000000000000) 
14'h01c2 : LOC =         127'b0000000000000000000001000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000200000008000000000000000000) 
14'h2f75 : LOC =         127'b0000000000000000000010000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000400000008000000000000000000) 
14'h316c : LOC =         127'b0000000000000000000100000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000800000008000000000000000000) 
14'h0d5e : LOC =         127'b0000000000000000001000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00001000000008000000000000000000) 
14'h364d : LOC =         127'b0000000000000000010000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00002000000008000000000000000000) 
14'h031c : LOC =         127'b0000000000000000100000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00004000000008000000000000000000) 
14'h2ac9 : LOC =         127'b0000000000000001000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00008000000008000000000000000000) 
14'h3a14 : LOC =         127'b0000000000000010000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00010000000008000000000000000000) 
14'h1bae : LOC =         127'b0000000000000100000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00020000000008000000000000000000) 
14'h1bad : LOC =         127'b0000000000001000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00040000000008000000000000000000) 
14'h1bab : LOC =         127'b0000000000010000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00080000000008000000000000000000) 
14'h1ba7 : LOC =         127'b0000000000100000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00100000000008000000000000000000) 
14'h1bbf : LOC =         127'b0000000001000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00200000000008000000000000000000) 
14'h1b8f : LOC =         127'b0000000010000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00400000000008000000000000000000) 
14'h1bef : LOC =         127'b0000000100000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00800000000008000000000000000000) 
14'h1b2f : LOC =         127'b0000001000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x01000000000008000000000000000000) 
14'h1aaf : LOC =         127'b0000010000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x02000000000008000000000000000000) 
14'h19af : LOC =         127'b0000100000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x04000000000008000000000000000000) 
14'h1faf : LOC =         127'b0001000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x08000000000008000000000000000000) 
14'h13af : LOC =         127'b0010000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x10000000000008000000000000000000) 
14'h0baf : LOC =         127'b0100000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x20000000000008000000000000000000) 
14'h3baf : LOC =         127'b1000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x40000000000008000000000000000000) 
14'h375e : LOC =         127'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000; // S (0x00000000000010000000000000000000) 
14'h1a95 : LOC =         127'b0000000000000000000000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000030000000000000000000) 
14'h2fbf : LOC =         127'b0000000000000000000000000000000000000000000000001010000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000050000000000000000000) 
14'h069c : LOC =         127'b0000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000090000000000000000000) 
14'h17ad : LOC =         127'b0000000000000000000000000000000000000000000000100010000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000110000000000000000000) 
14'h35cf : LOC =         127'b0000000000000000000000000000000000000000000001000010000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000210000000000000000000) 
14'h327c : LOC =         127'b0000000000000000000000000000000000000000000010000010000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000410000000000000000000) 
14'h3d1a : LOC =         127'b0000000000000000000000000000000000000000000100000010000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000810000000000000000000) 
14'h23d6 : LOC =         127'b0000000000000000000000000000000000000000001000000010000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000001010000000000000000000) 
14'h1e4e : LOC =         127'b0000000000000000000000000000000000000000010000000010000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000002010000000000000000000) 
14'h2609 : LOC =         127'b0000000000000000000000000000000000000000100000000010000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000004010000000000000000000) 
14'h15f0 : LOC =         127'b0000000000000000000000000000000000000001000000000010000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000008010000000000000000000) 
14'h3175 : LOC =         127'b0000000000000000000000000000000000000010000000000010000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000010010000000000000000000) 
14'h3b08 : LOC =         127'b0000000000000000000000000000000000000100000000000010000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000020010000000000000000000) 
14'h2ff2 : LOC =         127'b0000000000000000000000000000000000001000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000040010000000000000000000) 
14'h0606 : LOC =         127'b0000000000000000000000000000000000010000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000080010000000000000000000) 
14'h1699 : LOC =         127'b0000000000000000000000000000000000100000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000100010000000000000000000) 
14'h37a7 : LOC =         127'b0000000000000000000000000000000001000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000200010000000000000000000) 
14'h36ac : LOC =         127'b0000000000000000000000000000000010000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000400010000000000000000000) 
14'h34ba : LOC =         127'b0000000000000000000000000000000100000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000800010000000000000000000) 
14'h3096 : LOC =         127'b0000000000000000000000000000001000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000001000010000000000000000000) 
14'h38ce : LOC =         127'b0000000000000000000000000000010000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000002000010000000000000000000) 
14'h287e : LOC =         127'b0000000000000000000000000000100000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000004000010000000000000000000) 
14'h091e : LOC =         127'b0000000000000000000000000001000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000008000010000000000000000000) 
14'h08a9 : LOC =         127'b0000000000000000000000000010000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000010000010000000000000000000) 
14'h0bc7 : LOC =         127'b0000000000000000000000000100000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000020000010000000000000000000) 
14'h0d1b : LOC =         127'b0000000000000000000000001000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000040000010000000000000000000) 
14'h00a3 : LOC =         127'b0000000000000000000000010000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000080000010000000000000000000) 
14'h1bd3 : LOC =         127'b0000000000000000000000100000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000100000010000000000000000000) 
14'h2d33 : LOC =         127'b0000000000000000000001000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000200000010000000000000000000) 
14'h0384 : LOC =         127'b0000000000000000000010000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000400000010000000000000000000) 
14'h1d9d : LOC =         127'b0000000000000000000100000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000800000010000000000000000000) 
14'h21af : LOC =         127'b0000000000000000001000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00001000000010000000000000000000) 
14'h1abc : LOC =         127'b0000000000000000010000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00002000000010000000000000000000) 
14'h2fed : LOC =         127'b0000000000000000100000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00004000000010000000000000000000) 
14'h0638 : LOC =         127'b0000000000000001000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00008000000010000000000000000000) 
14'h16e5 : LOC =         127'b0000000000000010000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00010000000010000000000000000000) 
14'h375f : LOC =         127'b0000000000000100000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00020000000010000000000000000000) 
14'h375c : LOC =         127'b0000000000001000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00040000000010000000000000000000) 
14'h375a : LOC =         127'b0000000000010000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00080000000010000000000000000000) 
14'h3756 : LOC =         127'b0000000000100000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00100000000010000000000000000000) 
14'h374e : LOC =         127'b0000000001000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00200000000010000000000000000000) 
14'h377e : LOC =         127'b0000000010000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00400000000010000000000000000000) 
14'h371e : LOC =         127'b0000000100000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00800000000010000000000000000000) 
14'h37de : LOC =         127'b0000001000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x01000000000010000000000000000000) 
14'h365e : LOC =         127'b0000010000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x02000000000010000000000000000000) 
14'h355e : LOC =         127'b0000100000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x04000000000010000000000000000000) 
14'h335e : LOC =         127'b0001000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x08000000000010000000000000000000) 
14'h3f5e : LOC =         127'b0010000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x10000000000010000000000000000000) 
14'h275e : LOC =         127'b0100000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x20000000000010000000000000000000) 
14'h175e : LOC =         127'b1000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x40000000000010000000000000000000) 
14'h2dcb : LOC =         127'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000; // S (0x00000000000020000000000000000000) 
14'h352a : LOC =         127'b0000000000000000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000060000000000000000000) 
14'h1c09 : LOC =         127'b0000000000000000000000000000000000000000000000010100000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x000000000000a0000000000000000000) 
14'h0d38 : LOC =         127'b0000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000120000000000000000000) 
14'h2f5a : LOC =         127'b0000000000000000000000000000000000000000000001000100000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000220000000000000000000) 
14'h28e9 : LOC =         127'b0000000000000000000000000000000000000000000010000100000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000420000000000000000000) 
14'h278f : LOC =         127'b0000000000000000000000000000000000000000000100000100000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000820000000000000000000) 
14'h3943 : LOC =         127'b0000000000000000000000000000000000000000001000000100000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000001020000000000000000000) 
14'h04db : LOC =         127'b0000000000000000000000000000000000000000010000000100000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000002020000000000000000000) 
14'h3c9c : LOC =         127'b0000000000000000000000000000000000000000100000000100000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000004020000000000000000000) 
14'h0f65 : LOC =         127'b0000000000000000000000000000000000000001000000000100000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000008020000000000000000000) 
14'h2be0 : LOC =         127'b0000000000000000000000000000000000000010000000000100000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000010020000000000000000000) 
14'h219d : LOC =         127'b0000000000000000000000000000000000000100000000000100000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000020020000000000000000000) 
14'h3567 : LOC =         127'b0000000000000000000000000000000000001000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000040020000000000000000000) 
14'h1c93 : LOC =         127'b0000000000000000000000000000000000010000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000080020000000000000000000) 
14'h0c0c : LOC =         127'b0000000000000000000000000000000000100000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000100020000000000000000000) 
14'h2d32 : LOC =         127'b0000000000000000000000000000000001000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000200020000000000000000000) 
14'h2c39 : LOC =         127'b0000000000000000000000000000000010000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000400020000000000000000000) 
14'h2e2f : LOC =         127'b0000000000000000000000000000000100000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000800020000000000000000000) 
14'h2a03 : LOC =         127'b0000000000000000000000000000001000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000001000020000000000000000000) 
14'h225b : LOC =         127'b0000000000000000000000000000010000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000002000020000000000000000000) 
14'h32eb : LOC =         127'b0000000000000000000000000000100000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000004000020000000000000000000) 
14'h138b : LOC =         127'b0000000000000000000000000001000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000008000020000000000000000000) 
14'h123c : LOC =         127'b0000000000000000000000000010000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000010000020000000000000000000) 
14'h1152 : LOC =         127'b0000000000000000000000000100000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000020000020000000000000000000) 
14'h178e : LOC =         127'b0000000000000000000000001000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000040000020000000000000000000) 
14'h1a36 : LOC =         127'b0000000000000000000000010000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000080000020000000000000000000) 
14'h0146 : LOC =         127'b0000000000000000000000100000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000100000020000000000000000000) 
14'h37a6 : LOC =         127'b0000000000000000000001000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000200000020000000000000000000) 
14'h1911 : LOC =         127'b0000000000000000000010000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000400000020000000000000000000) 
14'h0708 : LOC =         127'b0000000000000000000100000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000800000020000000000000000000) 
14'h3b3a : LOC =         127'b0000000000000000001000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00001000000020000000000000000000) 
14'h0029 : LOC =         127'b0000000000000000010000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00002000000020000000000000000000) 
14'h3578 : LOC =         127'b0000000000000000100000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00004000000020000000000000000000) 
14'h1cad : LOC =         127'b0000000000000001000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00008000000020000000000000000000) 
14'h0c70 : LOC =         127'b0000000000000010000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00010000000020000000000000000000) 
14'h2dca : LOC =         127'b0000000000000100000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00020000000020000000000000000000) 
14'h2dc9 : LOC =         127'b0000000000001000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00040000000020000000000000000000) 
14'h2dcf : LOC =         127'b0000000000010000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00080000000020000000000000000000) 
14'h2dc3 : LOC =         127'b0000000000100000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00100000000020000000000000000000) 
14'h2ddb : LOC =         127'b0000000001000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00200000000020000000000000000000) 
14'h2deb : LOC =         127'b0000000010000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00400000000020000000000000000000) 
14'h2d8b : LOC =         127'b0000000100000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00800000000020000000000000000000) 
14'h2d4b : LOC =         127'b0000001000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x01000000000020000000000000000000) 
14'h2ccb : LOC =         127'b0000010000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x02000000000020000000000000000000) 
14'h2fcb : LOC =         127'b0000100000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x04000000000020000000000000000000) 
14'h29cb : LOC =         127'b0001000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x08000000000020000000000000000000) 
14'h25cb : LOC =         127'b0010000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x10000000000020000000000000000000) 
14'h3dcb : LOC =         127'b0100000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x20000000000020000000000000000000) 
14'h0dcb : LOC =         127'b1000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x40000000000020000000000000000000) 
14'h18e1 : LOC =         127'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000; // S (0x00000000000040000000000000000000) 
14'h2923 : LOC =         127'b0000000000000000000000000000000000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x000000000000c0000000000000000000) 
14'h3812 : LOC =         127'b0000000000000000000000000000000000000000000000101000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000140000000000000000000) 
14'h1a70 : LOC =         127'b0000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000240000000000000000000) 
14'h1dc3 : LOC =         127'b0000000000000000000000000000000000000000000010001000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000440000000000000000000) 
14'h12a5 : LOC =         127'b0000000000000000000000000000000000000000000100001000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000840000000000000000000) 
14'h0c69 : LOC =         127'b0000000000000000000000000000000000000000001000001000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000001040000000000000000000) 
14'h31f1 : LOC =         127'b0000000000000000000000000000000000000000010000001000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000002040000000000000000000) 
14'h09b6 : LOC =         127'b0000000000000000000000000000000000000000100000001000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000004040000000000000000000) 
14'h3a4f : LOC =         127'b0000000000000000000000000000000000000001000000001000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000008040000000000000000000) 
14'h1eca : LOC =         127'b0000000000000000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000010040000000000000000000) 
14'h14b7 : LOC =         127'b0000000000000000000000000000000000000100000000001000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000020040000000000000000000) 
14'h004d : LOC =         127'b0000000000000000000000000000000000001000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000040040000000000000000000) 
14'h29b9 : LOC =         127'b0000000000000000000000000000000000010000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000080040000000000000000000) 
14'h3926 : LOC =         127'b0000000000000000000000000000000000100000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000100040000000000000000000) 
14'h1818 : LOC =         127'b0000000000000000000000000000000001000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000200040000000000000000000) 
14'h1913 : LOC =         127'b0000000000000000000000000000000010000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000400040000000000000000000) 
14'h1b05 : LOC =         127'b0000000000000000000000000000000100000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000800040000000000000000000) 
14'h1f29 : LOC =         127'b0000000000000000000000000000001000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000001000040000000000000000000) 
14'h1771 : LOC =         127'b0000000000000000000000000000010000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000002000040000000000000000000) 
14'h07c1 : LOC =         127'b0000000000000000000000000000100000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000004000040000000000000000000) 
14'h26a1 : LOC =         127'b0000000000000000000000000001000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000008000040000000000000000000) 
14'h2716 : LOC =         127'b0000000000000000000000000010000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000010000040000000000000000000) 
14'h2478 : LOC =         127'b0000000000000000000000000100000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000020000040000000000000000000) 
14'h22a4 : LOC =         127'b0000000000000000000000001000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000040000040000000000000000000) 
14'h2f1c : LOC =         127'b0000000000000000000000010000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000080000040000000000000000000) 
14'h346c : LOC =         127'b0000000000000000000000100000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000100000040000000000000000000) 
14'h028c : LOC =         127'b0000000000000000000001000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000200000040000000000000000000) 
14'h2c3b : LOC =         127'b0000000000000000000010000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000400000040000000000000000000) 
14'h3222 : LOC =         127'b0000000000000000000100000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000800000040000000000000000000) 
14'h0e10 : LOC =         127'b0000000000000000001000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00001000000040000000000000000000) 
14'h3503 : LOC =         127'b0000000000000000010000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00002000000040000000000000000000) 
14'h0052 : LOC =         127'b0000000000000000100000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00004000000040000000000000000000) 
14'h2987 : LOC =         127'b0000000000000001000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00008000000040000000000000000000) 
14'h395a : LOC =         127'b0000000000000010000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00010000000040000000000000000000) 
14'h18e0 : LOC =         127'b0000000000000100000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00020000000040000000000000000000) 
14'h18e3 : LOC =         127'b0000000000001000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00040000000040000000000000000000) 
14'h18e5 : LOC =         127'b0000000000010000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00080000000040000000000000000000) 
14'h18e9 : LOC =         127'b0000000000100000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00100000000040000000000000000000) 
14'h18f1 : LOC =         127'b0000000001000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00200000000040000000000000000000) 
14'h18c1 : LOC =         127'b0000000010000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00400000000040000000000000000000) 
14'h18a1 : LOC =         127'b0000000100000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00800000000040000000000000000000) 
14'h1861 : LOC =         127'b0000001000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x01000000000040000000000000000000) 
14'h19e1 : LOC =         127'b0000010000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x02000000000040000000000000000000) 
14'h1ae1 : LOC =         127'b0000100000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x04000000000040000000000000000000) 
14'h1ce1 : LOC =         127'b0001000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x08000000000040000000000000000000) 
14'h10e1 : LOC =         127'b0010000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x10000000000040000000000000000000) 
14'h08e1 : LOC =         127'b0100000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x20000000000040000000000000000000) 
14'h38e1 : LOC =         127'b1000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x40000000000040000000000000000000) 
14'h31c2 : LOC =         127'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000; // S (0x00000000000080000000000000000000) 
14'h1131 : LOC =         127'b0000000000000000000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000180000000000000000000) 
14'h3353 : LOC =         127'b0000000000000000000000000000000000000000000001010000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000280000000000000000000) 
14'h34e0 : LOC =         127'b0000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000480000000000000000000) 
14'h3b86 : LOC =         127'b0000000000000000000000000000000000000000000100010000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000880000000000000000000) 
14'h254a : LOC =         127'b0000000000000000000000000000000000000000001000010000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000001080000000000000000000) 
14'h18d2 : LOC =         127'b0000000000000000000000000000000000000000010000010000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000002080000000000000000000) 
14'h2095 : LOC =         127'b0000000000000000000000000000000000000000100000010000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000004080000000000000000000) 
14'h136c : LOC =         127'b0000000000000000000000000000000000000001000000010000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000008080000000000000000000) 
14'h37e9 : LOC =         127'b0000000000000000000000000000000000000010000000010000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000010080000000000000000000) 
14'h3d94 : LOC =         127'b0000000000000000000000000000000000000100000000010000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000020080000000000000000000) 
14'h296e : LOC =         127'b0000000000000000000000000000000000001000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000040080000000000000000000) 
14'h009a : LOC =         127'b0000000000000000000000000000000000010000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000080080000000000000000000) 
14'h1005 : LOC =         127'b0000000000000000000000000000000000100000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000100080000000000000000000) 
14'h313b : LOC =         127'b0000000000000000000000000000000001000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000200080000000000000000000) 
14'h3030 : LOC =         127'b0000000000000000000000000000000010000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000400080000000000000000000) 
14'h3226 : LOC =         127'b0000000000000000000000000000000100000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000800080000000000000000000) 
14'h360a : LOC =         127'b0000000000000000000000000000001000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000001000080000000000000000000) 
14'h3e52 : LOC =         127'b0000000000000000000000000000010000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000002000080000000000000000000) 
14'h2ee2 : LOC =         127'b0000000000000000000000000000100000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000004000080000000000000000000) 
14'h0f82 : LOC =         127'b0000000000000000000000000001000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000008000080000000000000000000) 
14'h0e35 : LOC =         127'b0000000000000000000000000010000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000010000080000000000000000000) 
14'h0d5b : LOC =         127'b0000000000000000000000000100000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000020000080000000000000000000) 
14'h0b87 : LOC =         127'b0000000000000000000000001000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000040000080000000000000000000) 
14'h063f : LOC =         127'b0000000000000000000000010000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000080000080000000000000000000) 
14'h1d4f : LOC =         127'b0000000000000000000000100000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000100000080000000000000000000) 
14'h2baf : LOC =         127'b0000000000000000000001000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000200000080000000000000000000) 
14'h0518 : LOC =         127'b0000000000000000000010000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000400000080000000000000000000) 
14'h1b01 : LOC =         127'b0000000000000000000100000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000800000080000000000000000000) 
14'h2733 : LOC =         127'b0000000000000000001000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00001000000080000000000000000000) 
14'h1c20 : LOC =         127'b0000000000000000010000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00002000000080000000000000000000) 
14'h2971 : LOC =         127'b0000000000000000100000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00004000000080000000000000000000) 
14'h00a4 : LOC =         127'b0000000000000001000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00008000000080000000000000000000) 
14'h1079 : LOC =         127'b0000000000000010000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00010000000080000000000000000000) 
14'h31c3 : LOC =         127'b0000000000000100000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00020000000080000000000000000000) 
14'h31c0 : LOC =         127'b0000000000001000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00040000000080000000000000000000) 
14'h31c6 : LOC =         127'b0000000000010000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00080000000080000000000000000000) 
14'h31ca : LOC =         127'b0000000000100000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00100000000080000000000000000000) 
14'h31d2 : LOC =         127'b0000000001000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00200000000080000000000000000000) 
14'h31e2 : LOC =         127'b0000000010000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00400000000080000000000000000000) 
14'h3182 : LOC =         127'b0000000100000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00800000000080000000000000000000) 
14'h3142 : LOC =         127'b0000001000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x01000000000080000000000000000000) 
14'h30c2 : LOC =         127'b0000010000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x02000000000080000000000000000000) 
14'h33c2 : LOC =         127'b0000100000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x04000000000080000000000000000000) 
14'h35c2 : LOC =         127'b0001000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x08000000000080000000000000000000) 
14'h39c2 : LOC =         127'b0010000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x10000000000080000000000000000000) 
14'h21c2 : LOC =         127'b0100000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x20000000000080000000000000000000) 
14'h11c2 : LOC =         127'b1000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x40000000000080000000000000000000) 
14'h20f3 : LOC =         127'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000; // S (0x00000000000100000000000000000000) 
14'h2262 : LOC =         127'b0000000000000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000300000000000000000000) 
14'h25d1 : LOC =         127'b0000000000000000000000000000000000000000000010100000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000500000000000000000000) 
14'h2ab7 : LOC =         127'b0000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000900000000000000000000) 
14'h347b : LOC =         127'b0000000000000000000000000000000000000000001000100000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000001100000000000000000000) 
14'h09e3 : LOC =         127'b0000000000000000000000000000000000000000010000100000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000002100000000000000000000) 
14'h31a4 : LOC =         127'b0000000000000000000000000000000000000000100000100000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000004100000000000000000000) 
14'h025d : LOC =         127'b0000000000000000000000000000000000000001000000100000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000008100000000000000000000) 
14'h26d8 : LOC =         127'b0000000000000000000000000000000000000010000000100000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000010100000000000000000000) 
14'h2ca5 : LOC =         127'b0000000000000000000000000000000000000100000000100000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000020100000000000000000000) 
14'h385f : LOC =         127'b0000000000000000000000000000000000001000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000040100000000000000000000) 
14'h11ab : LOC =         127'b0000000000000000000000000000000000010000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000080100000000000000000000) 
14'h0134 : LOC =         127'b0000000000000000000000000000000000100000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000100100000000000000000000) 
14'h200a : LOC =         127'b0000000000000000000000000000000001000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000200100000000000000000000) 
14'h2101 : LOC =         127'b0000000000000000000000000000000010000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000400100000000000000000000) 
14'h2317 : LOC =         127'b0000000000000000000000000000000100000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000800100000000000000000000) 
14'h273b : LOC =         127'b0000000000000000000000000000001000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000001000100000000000000000000) 
14'h2f63 : LOC =         127'b0000000000000000000000000000010000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000002000100000000000000000000) 
14'h3fd3 : LOC =         127'b0000000000000000000000000000100000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000004000100000000000000000000) 
14'h1eb3 : LOC =         127'b0000000000000000000000000001000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000008000100000000000000000000) 
14'h1f04 : LOC =         127'b0000000000000000000000000010000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000010000100000000000000000000) 
14'h1c6a : LOC =         127'b0000000000000000000000000100000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000020000100000000000000000000) 
14'h1ab6 : LOC =         127'b0000000000000000000000001000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000040000100000000000000000000) 
14'h170e : LOC =         127'b0000000000000000000000010000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000080000100000000000000000000) 
14'h0c7e : LOC =         127'b0000000000000000000000100000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000100000100000000000000000000) 
14'h3a9e : LOC =         127'b0000000000000000000001000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000200000100000000000000000000) 
14'h1429 : LOC =         127'b0000000000000000000010000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000400000100000000000000000000) 
14'h0a30 : LOC =         127'b0000000000000000000100000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000800000100000000000000000000) 
14'h3602 : LOC =         127'b0000000000000000001000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00001000000100000000000000000000) 
14'h0d11 : LOC =         127'b0000000000000000010000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00002000000100000000000000000000) 
14'h3840 : LOC =         127'b0000000000000000100000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00004000000100000000000000000000) 
14'h1195 : LOC =         127'b0000000000000001000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00008000000100000000000000000000) 
14'h0148 : LOC =         127'b0000000000000010000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00010000000100000000000000000000) 
14'h20f2 : LOC =         127'b0000000000000100000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00020000000100000000000000000000) 
14'h20f1 : LOC =         127'b0000000000001000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00040000000100000000000000000000) 
14'h20f7 : LOC =         127'b0000000000010000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00080000000100000000000000000000) 
14'h20fb : LOC =         127'b0000000000100000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00100000000100000000000000000000) 
14'h20e3 : LOC =         127'b0000000001000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00200000000100000000000000000000) 
14'h20d3 : LOC =         127'b0000000010000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00400000000100000000000000000000) 
14'h20b3 : LOC =         127'b0000000100000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00800000000100000000000000000000) 
14'h2073 : LOC =         127'b0000001000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x01000000000100000000000000000000) 
14'h21f3 : LOC =         127'b0000010000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x02000000000100000000000000000000) 
14'h22f3 : LOC =         127'b0000100000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x04000000000100000000000000000000) 
14'h24f3 : LOC =         127'b0001000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x08000000000100000000000000000000) 
14'h28f3 : LOC =         127'b0010000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x10000000000100000000000000000000) 
14'h30f3 : LOC =         127'b0100000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x20000000000100000000000000000000) 
14'h00f3 : LOC =         127'b1000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x40000000000100000000000000000000) 
14'h0291 : LOC =         127'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000; // S (0x00000000000200000000000000000000) 
14'h07b3 : LOC =         127'b0000000000000000000000000000000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000600000000000000000000) 
14'h08d5 : LOC =         127'b0000000000000000000000000000000000000000000101000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000a00000000000000000000) 
14'h1619 : LOC =         127'b0000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000001200000000000000000000) 
14'h2b81 : LOC =         127'b0000000000000000000000000000000000000000010001000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000002200000000000000000000) 
14'h13c6 : LOC =         127'b0000000000000000000000000000000000000000100001000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000004200000000000000000000) 
14'h203f : LOC =         127'b0000000000000000000000000000000000000001000001000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000008200000000000000000000) 
14'h04ba : LOC =         127'b0000000000000000000000000000000000000010000001000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000010200000000000000000000) 
14'h0ec7 : LOC =         127'b0000000000000000000000000000000000000100000001000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000020200000000000000000000) 
14'h1a3d : LOC =         127'b0000000000000000000000000000000000001000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000040200000000000000000000) 
14'h33c9 : LOC =         127'b0000000000000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000080200000000000000000000) 
14'h2356 : LOC =         127'b0000000000000000000000000000000000100000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000100200000000000000000000) 
14'h0268 : LOC =         127'b0000000000000000000000000000000001000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000200200000000000000000000) 
14'h0363 : LOC =         127'b0000000000000000000000000000000010000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000400200000000000000000000) 
14'h0175 : LOC =         127'b0000000000000000000000000000000100000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000800200000000000000000000) 
14'h0559 : LOC =         127'b0000000000000000000000000000001000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000001000200000000000000000000) 
14'h0d01 : LOC =         127'b0000000000000000000000000000010000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000002000200000000000000000000) 
14'h1db1 : LOC =         127'b0000000000000000000000000000100000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000004000200000000000000000000) 
14'h3cd1 : LOC =         127'b0000000000000000000000000001000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000008000200000000000000000000) 
14'h3d66 : LOC =         127'b0000000000000000000000000010000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000010000200000000000000000000) 
14'h3e08 : LOC =         127'b0000000000000000000000000100000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000020000200000000000000000000) 
14'h38d4 : LOC =         127'b0000000000000000000000001000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000040000200000000000000000000) 
14'h356c : LOC =         127'b0000000000000000000000010000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000080000200000000000000000000) 
14'h2e1c : LOC =         127'b0000000000000000000000100000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000100000200000000000000000000) 
14'h18fc : LOC =         127'b0000000000000000000001000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000200000200000000000000000000) 
14'h364b : LOC =         127'b0000000000000000000010000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000400000200000000000000000000) 
14'h2852 : LOC =         127'b0000000000000000000100000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000800000200000000000000000000) 
14'h1460 : LOC =         127'b0000000000000000001000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00001000000200000000000000000000) 
14'h2f73 : LOC =         127'b0000000000000000010000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00002000000200000000000000000000) 
14'h1a22 : LOC =         127'b0000000000000000100000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00004000000200000000000000000000) 
14'h33f7 : LOC =         127'b0000000000000001000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00008000000200000000000000000000) 
14'h232a : LOC =         127'b0000000000000010000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00010000000200000000000000000000) 
14'h0290 : LOC =         127'b0000000000000100000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00020000000200000000000000000000) 
14'h0293 : LOC =         127'b0000000000001000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00040000000200000000000000000000) 
14'h0295 : LOC =         127'b0000000000010000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00080000000200000000000000000000) 
14'h0299 : LOC =         127'b0000000000100000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00100000000200000000000000000000) 
14'h0281 : LOC =         127'b0000000001000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00200000000200000000000000000000) 
14'h02b1 : LOC =         127'b0000000010000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00400000000200000000000000000000) 
14'h02d1 : LOC =         127'b0000000100000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00800000000200000000000000000000) 
14'h0211 : LOC =         127'b0000001000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x01000000000200000000000000000000) 
14'h0391 : LOC =         127'b0000010000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x02000000000200000000000000000000) 
14'h0091 : LOC =         127'b0000100000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x04000000000200000000000000000000) 
14'h0691 : LOC =         127'b0001000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x08000000000200000000000000000000) 
14'h0a91 : LOC =         127'b0010000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x10000000000200000000000000000000) 
14'h1291 : LOC =         127'b0100000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x20000000000200000000000000000000) 
14'h2291 : LOC =         127'b1000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x40000000000200000000000000000000) 
14'h0522 : LOC =         127'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000; // S (0x00000000000400000000000000000000) 
14'h0f66 : LOC =         127'b0000000000000000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000000c00000000000000000000) 
14'h11aa : LOC =         127'b0000000000000000000000000000000000000000001010000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000001400000000000000000000) 
14'h2c32 : LOC =         127'b0000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000002400000000000000000000) 
14'h1475 : LOC =         127'b0000000000000000000000000000000000000000100010000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000004400000000000000000000) 
14'h278c : LOC =         127'b0000000000000000000000000000000000000001000010000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000008400000000000000000000) 
14'h0309 : LOC =         127'b0000000000000000000000000000000000000010000010000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000010400000000000000000000) 
14'h0974 : LOC =         127'b0000000000000000000000000000000000000100000010000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000020400000000000000000000) 
14'h1d8e : LOC =         127'b0000000000000000000000000000000000001000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000040400000000000000000000) 
14'h347a : LOC =         127'b0000000000000000000000000000000000010000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000080400000000000000000000) 
14'h24e5 : LOC =         127'b0000000000000000000000000000000000100000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000100400000000000000000000) 
14'h05db : LOC =         127'b0000000000000000000000000000000001000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000200400000000000000000000) 
14'h04d0 : LOC =         127'b0000000000000000000000000000000010000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000400400000000000000000000) 
14'h06c6 : LOC =         127'b0000000000000000000000000000000100000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000800400000000000000000000) 
14'h02ea : LOC =         127'b0000000000000000000000000000001000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000001000400000000000000000000) 
14'h0ab2 : LOC =         127'b0000000000000000000000000000010000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000002000400000000000000000000) 
14'h1a02 : LOC =         127'b0000000000000000000000000000100000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000004000400000000000000000000) 
14'h3b62 : LOC =         127'b0000000000000000000000000001000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000008000400000000000000000000) 
14'h3ad5 : LOC =         127'b0000000000000000000000000010000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000010000400000000000000000000) 
14'h39bb : LOC =         127'b0000000000000000000000000100000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000020000400000000000000000000) 
14'h3f67 : LOC =         127'b0000000000000000000000001000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000040000400000000000000000000) 
14'h32df : LOC =         127'b0000000000000000000000010000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000080000400000000000000000000) 
14'h29af : LOC =         127'b0000000000000000000000100000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000100000400000000000000000000) 
14'h1f4f : LOC =         127'b0000000000000000000001000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000200000400000000000000000000) 
14'h31f8 : LOC =         127'b0000000000000000000010000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000400000400000000000000000000) 
14'h2fe1 : LOC =         127'b0000000000000000000100000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000800000400000000000000000000) 
14'h13d3 : LOC =         127'b0000000000000000001000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00001000000400000000000000000000) 
14'h28c0 : LOC =         127'b0000000000000000010000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00002000000400000000000000000000) 
14'h1d91 : LOC =         127'b0000000000000000100000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00004000000400000000000000000000) 
14'h3444 : LOC =         127'b0000000000000001000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00008000000400000000000000000000) 
14'h2499 : LOC =         127'b0000000000000010000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00010000000400000000000000000000) 
14'h0523 : LOC =         127'b0000000000000100000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00020000000400000000000000000000) 
14'h0520 : LOC =         127'b0000000000001000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00040000000400000000000000000000) 
14'h0526 : LOC =         127'b0000000000010000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00080000000400000000000000000000) 
14'h052a : LOC =         127'b0000000000100000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00100000000400000000000000000000) 
14'h0532 : LOC =         127'b0000000001000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00200000000400000000000000000000) 
14'h0502 : LOC =         127'b0000000010000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00400000000400000000000000000000) 
14'h0562 : LOC =         127'b0000000100000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00800000000400000000000000000000) 
14'h05a2 : LOC =         127'b0000001000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x01000000000400000000000000000000) 
14'h0422 : LOC =         127'b0000010000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x02000000000400000000000000000000) 
14'h0722 : LOC =         127'b0000100000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x04000000000400000000000000000000) 
14'h0122 : LOC =         127'b0001000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x08000000000400000000000000000000) 
14'h0d22 : LOC =         127'b0010000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x10000000000400000000000000000000) 
14'h1522 : LOC =         127'b0100000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x20000000000400000000000000000000) 
14'h2522 : LOC =         127'b1000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x40000000000400000000000000000000) 
14'h0a44 : LOC =         127'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000; // S (0x00000000000800000000000000000000) 
14'h1ecc : LOC =         127'b0000000000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000001800000000000000000000) 
14'h2354 : LOC =         127'b0000000000000000000000000000000000000000010100000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000002800000000000000000000) 
14'h1b13 : LOC =         127'b0000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000004800000000000000000000) 
14'h28ea : LOC =         127'b0000000000000000000000000000000000000001000100000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000008800000000000000000000) 
14'h0c6f : LOC =         127'b0000000000000000000000000000000000000010000100000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000010800000000000000000000) 
14'h0612 : LOC =         127'b0000000000000000000000000000000000000100000100000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000020800000000000000000000) 
14'h12e8 : LOC =         127'b0000000000000000000000000000000000001000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000040800000000000000000000) 
14'h3b1c : LOC =         127'b0000000000000000000000000000000000010000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000080800000000000000000000) 
14'h2b83 : LOC =         127'b0000000000000000000000000000000000100000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000100800000000000000000000) 
14'h0abd : LOC =         127'b0000000000000000000000000000000001000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000200800000000000000000000) 
14'h0bb6 : LOC =         127'b0000000000000000000000000000000010000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000400800000000000000000000) 
14'h09a0 : LOC =         127'b0000000000000000000000000000000100000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000800800000000000000000000) 
14'h0d8c : LOC =         127'b0000000000000000000000000000001000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000001000800000000000000000000) 
14'h05d4 : LOC =         127'b0000000000000000000000000000010000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000002000800000000000000000000) 
14'h1564 : LOC =         127'b0000000000000000000000000000100000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000004000800000000000000000000) 
14'h3404 : LOC =         127'b0000000000000000000000000001000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000008000800000000000000000000) 
14'h35b3 : LOC =         127'b0000000000000000000000000010000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000010000800000000000000000000) 
14'h36dd : LOC =         127'b0000000000000000000000000100000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000020000800000000000000000000) 
14'h3001 : LOC =         127'b0000000000000000000000001000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000040000800000000000000000000) 
14'h3db9 : LOC =         127'b0000000000000000000000010000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000080000800000000000000000000) 
14'h26c9 : LOC =         127'b0000000000000000000000100000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000100000800000000000000000000) 
14'h1029 : LOC =         127'b0000000000000000000001000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000200000800000000000000000000) 
14'h3e9e : LOC =         127'b0000000000000000000010000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000400000800000000000000000000) 
14'h2087 : LOC =         127'b0000000000000000000100000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000800000800000000000000000000) 
14'h1cb5 : LOC =         127'b0000000000000000001000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00001000000800000000000000000000) 
14'h27a6 : LOC =         127'b0000000000000000010000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00002000000800000000000000000000) 
14'h12f7 : LOC =         127'b0000000000000000100000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00004000000800000000000000000000) 
14'h3b22 : LOC =         127'b0000000000000001000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00008000000800000000000000000000) 
14'h2bff : LOC =         127'b0000000000000010000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00010000000800000000000000000000) 
14'h0a45 : LOC =         127'b0000000000000100000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00020000000800000000000000000000) 
14'h0a46 : LOC =         127'b0000000000001000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00040000000800000000000000000000) 
14'h0a40 : LOC =         127'b0000000000010000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00080000000800000000000000000000) 
14'h0a4c : LOC =         127'b0000000000100000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00100000000800000000000000000000) 
14'h0a54 : LOC =         127'b0000000001000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00200000000800000000000000000000) 
14'h0a64 : LOC =         127'b0000000010000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00400000000800000000000000000000) 
14'h0a04 : LOC =         127'b0000000100000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00800000000800000000000000000000) 
14'h0ac4 : LOC =         127'b0000001000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x01000000000800000000000000000000) 
14'h0b44 : LOC =         127'b0000010000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x02000000000800000000000000000000) 
14'h0844 : LOC =         127'b0000100000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x04000000000800000000000000000000) 
14'h0e44 : LOC =         127'b0001000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x08000000000800000000000000000000) 
14'h0244 : LOC =         127'b0010000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x10000000000800000000000000000000) 
14'h1a44 : LOC =         127'b0100000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x20000000000800000000000000000000) 
14'h2a44 : LOC =         127'b1000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x40000000000800000000000000000000) 
14'h1488 : LOC =         127'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // S (0x00000000001000000000000000000000) 
14'h3d98 : LOC =         127'b0000000000000000000000000000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000003000000000000000000000) 
14'h05df : LOC =         127'b0000000000000000000000000000000000000000101000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000005000000000000000000000) 
14'h3626 : LOC =         127'b0000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000009000000000000000000000) 
14'h12a3 : LOC =         127'b0000000000000000000000000000000000000010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000011000000000000000000000) 
14'h18de : LOC =         127'b0000000000000000000000000000000000000100001000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000021000000000000000000000) 
14'h0c24 : LOC =         127'b0000000000000000000000000000000000001000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000041000000000000000000000) 
14'h25d0 : LOC =         127'b0000000000000000000000000000000000010000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000081000000000000000000000) 
14'h354f : LOC =         127'b0000000000000000000000000000000000100000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000101000000000000000000000) 
14'h1471 : LOC =         127'b0000000000000000000000000000000001000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000201000000000000000000000) 
14'h157a : LOC =         127'b0000000000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000401000000000000000000000) 
14'h176c : LOC =         127'b0000000000000000000000000000000100000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000801000000000000000000000) 
14'h1340 : LOC =         127'b0000000000000000000000000000001000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000001001000000000000000000000) 
14'h1b18 : LOC =         127'b0000000000000000000000000000010000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000002001000000000000000000000) 
14'h0ba8 : LOC =         127'b0000000000000000000000000000100000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000004001000000000000000000000) 
14'h2ac8 : LOC =         127'b0000000000000000000000000001000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000008001000000000000000000000) 
14'h2b7f : LOC =         127'b0000000000000000000000000010000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000010001000000000000000000000) 
14'h2811 : LOC =         127'b0000000000000000000000000100000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000020001000000000000000000000) 
14'h2ecd : LOC =         127'b0000000000000000000000001000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000040001000000000000000000000) 
14'h2375 : LOC =         127'b0000000000000000000000010000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000080001000000000000000000000) 
14'h3805 : LOC =         127'b0000000000000000000000100000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000100001000000000000000000000) 
14'h0ee5 : LOC =         127'b0000000000000000000001000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000200001000000000000000000000) 
14'h2052 : LOC =         127'b0000000000000000000010000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000400001000000000000000000000) 
14'h3e4b : LOC =         127'b0000000000000000000100000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000800001000000000000000000000) 
14'h0279 : LOC =         127'b0000000000000000001000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00001000001000000000000000000000) 
14'h396a : LOC =         127'b0000000000000000010000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00002000001000000000000000000000) 
14'h0c3b : LOC =         127'b0000000000000000100000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00004000001000000000000000000000) 
14'h25ee : LOC =         127'b0000000000000001000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00008000001000000000000000000000) 
14'h3533 : LOC =         127'b0000000000000010000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00010000001000000000000000000000) 
14'h1489 : LOC =         127'b0000000000000100000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00020000001000000000000000000000) 
14'h148a : LOC =         127'b0000000000001000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00040000001000000000000000000000) 
14'h148c : LOC =         127'b0000000000010000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00080000001000000000000000000000) 
14'h1480 : LOC =         127'b0000000000100000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00100000001000000000000000000000) 
14'h1498 : LOC =         127'b0000000001000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00200000001000000000000000000000) 
14'h14a8 : LOC =         127'b0000000010000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00400000001000000000000000000000) 
14'h14c8 : LOC =         127'b0000000100000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00800000001000000000000000000000) 
14'h1408 : LOC =         127'b0000001000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x01000000001000000000000000000000) 
14'h1588 : LOC =         127'b0000010000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x02000000001000000000000000000000) 
14'h1688 : LOC =         127'b0000100000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x04000000001000000000000000000000) 
14'h1088 : LOC =         127'b0001000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x08000000001000000000000000000000) 
14'h1c88 : LOC =         127'b0010000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x10000000001000000000000000000000) 
14'h0488 : LOC =         127'b0100000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x20000000001000000000000000000000) 
14'h3488 : LOC =         127'b1000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x40000000001000000000000000000000) 
14'h2910 : LOC =         127'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // S (0x00000000002000000000000000000000) 
14'h3847 : LOC =         127'b0000000000000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000006000000000000000000000) 
14'h0bbe : LOC =         127'b0000000000000000000000000000000000000001010000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x0000000000a000000000000000000000) 
14'h2f3b : LOC =         127'b0000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000012000000000000000000000) 
14'h2546 : LOC =         127'b0000000000000000000000000000000000000100010000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000022000000000000000000000) 
14'h31bc : LOC =         127'b0000000000000000000000000000000000001000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000042000000000000000000000) 
14'h1848 : LOC =         127'b0000000000000000000000000000000000010000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000082000000000000000000000) 
14'h08d7 : LOC =         127'b0000000000000000000000000000000000100000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000102000000000000000000000) 
14'h29e9 : LOC =         127'b0000000000000000000000000000000001000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000202000000000000000000000) 
14'h28e2 : LOC =         127'b0000000000000000000000000000000010000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000402000000000000000000000) 
14'h2af4 : LOC =         127'b0000000000000000000000000000000100000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000802000000000000000000000) 
14'h2ed8 : LOC =         127'b0000000000000000000000000000001000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000001002000000000000000000000) 
14'h2680 : LOC =         127'b0000000000000000000000000000010000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000002002000000000000000000000) 
14'h3630 : LOC =         127'b0000000000000000000000000000100000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000004002000000000000000000000) 
14'h1750 : LOC =         127'b0000000000000000000000000001000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000008002000000000000000000000) 
14'h16e7 : LOC =         127'b0000000000000000000000000010000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000010002000000000000000000000) 
14'h1589 : LOC =         127'b0000000000000000000000000100000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000020002000000000000000000000) 
14'h1355 : LOC =         127'b0000000000000000000000001000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000040002000000000000000000000) 
14'h1eed : LOC =         127'b0000000000000000000000010000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000080002000000000000000000000) 
14'h059d : LOC =         127'b0000000000000000000000100000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000100002000000000000000000000) 
14'h337d : LOC =         127'b0000000000000000000001000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000200002000000000000000000000) 
14'h1dca : LOC =         127'b0000000000000000000010000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000400002000000000000000000000) 
14'h03d3 : LOC =         127'b0000000000000000000100000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000800002000000000000000000000) 
14'h3fe1 : LOC =         127'b0000000000000000001000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00001000002000000000000000000000) 
14'h04f2 : LOC =         127'b0000000000000000010000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00002000002000000000000000000000) 
14'h31a3 : LOC =         127'b0000000000000000100000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00004000002000000000000000000000) 
14'h1876 : LOC =         127'b0000000000000001000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00008000002000000000000000000000) 
14'h08ab : LOC =         127'b0000000000000010000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00010000002000000000000000000000) 
14'h2911 : LOC =         127'b0000000000000100000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00020000002000000000000000000000) 
14'h2912 : LOC =         127'b0000000000001000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00040000002000000000000000000000) 
14'h2914 : LOC =         127'b0000000000010000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00080000002000000000000000000000) 
14'h2918 : LOC =         127'b0000000000100000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00100000002000000000000000000000) 
14'h2900 : LOC =         127'b0000000001000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00200000002000000000000000000000) 
14'h2930 : LOC =         127'b0000000010000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00400000002000000000000000000000) 
14'h2950 : LOC =         127'b0000000100000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00800000002000000000000000000000) 
14'h2990 : LOC =         127'b0000001000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x01000000002000000000000000000000) 
14'h2810 : LOC =         127'b0000010000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x02000000002000000000000000000000) 
14'h2b10 : LOC =         127'b0000100000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x04000000002000000000000000000000) 
14'h2d10 : LOC =         127'b0001000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x08000000002000000000000000000000) 
14'h2110 : LOC =         127'b0010000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x10000000002000000000000000000000) 
14'h3910 : LOC =         127'b0100000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x20000000002000000000000000000000) 
14'h0910 : LOC =         127'b1000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x40000000002000000000000000000000) 
14'h1157 : LOC =         127'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // S (0x00000000004000000000000000000000) 
14'h33f9 : LOC =         127'b0000000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x0000000000c000000000000000000000) 
14'h177c : LOC =         127'b0000000000000000000000000000000000000010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000014000000000000000000000) 
14'h1d01 : LOC =         127'b0000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000024000000000000000000000) 
14'h09fb : LOC =         127'b0000000000000000000000000000000000001000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000044000000000000000000000) 
14'h200f : LOC =         127'b0000000000000000000000000000000000010000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000084000000000000000000000) 
14'h3090 : LOC =         127'b0000000000000000000000000000000000100000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000104000000000000000000000) 
14'h11ae : LOC =         127'b0000000000000000000000000000000001000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000204000000000000000000000) 
14'h10a5 : LOC =         127'b0000000000000000000000000000000010000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000404000000000000000000000) 
14'h12b3 : LOC =         127'b0000000000000000000000000000000100000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000804000000000000000000000) 
14'h169f : LOC =         127'b0000000000000000000000000000001000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000001004000000000000000000000) 
14'h1ec7 : LOC =         127'b0000000000000000000000000000010000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000002004000000000000000000000) 
14'h0e77 : LOC =         127'b0000000000000000000000000000100000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000004004000000000000000000000) 
14'h2f17 : LOC =         127'b0000000000000000000000000001000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000008004000000000000000000000) 
14'h2ea0 : LOC =         127'b0000000000000000000000000010000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000010004000000000000000000000) 
14'h2dce : LOC =         127'b0000000000000000000000000100000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000020004000000000000000000000) 
14'h2b12 : LOC =         127'b0000000000000000000000001000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000040004000000000000000000000) 
14'h26aa : LOC =         127'b0000000000000000000000010000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000080004000000000000000000000) 
14'h3dda : LOC =         127'b0000000000000000000000100000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000100004000000000000000000000) 
14'h0b3a : LOC =         127'b0000000000000000000001000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000200004000000000000000000000) 
14'h258d : LOC =         127'b0000000000000000000010000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000400004000000000000000000000) 
14'h3b94 : LOC =         127'b0000000000000000000100000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000800004000000000000000000000) 
14'h07a6 : LOC =         127'b0000000000000000001000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00001000004000000000000000000000) 
14'h3cb5 : LOC =         127'b0000000000000000010000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00002000004000000000000000000000) 
14'h09e4 : LOC =         127'b0000000000000000100000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00004000004000000000000000000000) 
14'h2031 : LOC =         127'b0000000000000001000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00008000004000000000000000000000) 
14'h30ec : LOC =         127'b0000000000000010000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00010000004000000000000000000000) 
14'h1156 : LOC =         127'b0000000000000100000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00020000004000000000000000000000) 
14'h1155 : LOC =         127'b0000000000001000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00040000004000000000000000000000) 
14'h1153 : LOC =         127'b0000000000010000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00080000004000000000000000000000) 
14'h115f : LOC =         127'b0000000000100000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00100000004000000000000000000000) 
14'h1147 : LOC =         127'b0000000001000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00200000004000000000000000000000) 
14'h1177 : LOC =         127'b0000000010000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00400000004000000000000000000000) 
14'h1117 : LOC =         127'b0000000100000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00800000004000000000000000000000) 
14'h11d7 : LOC =         127'b0000001000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x01000000004000000000000000000000) 
14'h1057 : LOC =         127'b0000010000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x02000000004000000000000000000000) 
14'h1357 : LOC =         127'b0000100000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x04000000004000000000000000000000) 
14'h1557 : LOC =         127'b0001000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x08000000004000000000000000000000) 
14'h1957 : LOC =         127'b0010000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x10000000004000000000000000000000) 
14'h0157 : LOC =         127'b0100000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x20000000004000000000000000000000) 
14'h3157 : LOC =         127'b1000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x40000000004000000000000000000000) 
14'h22ae : LOC =         127'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // S (0x00000000008000000000000000000000) 
14'h2485 : LOC =         127'b0000000000000000000000000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000018000000000000000000000) 
14'h2ef8 : LOC =         127'b0000000000000000000000000000000000000101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000028000000000000000000000) 
14'h3a02 : LOC =         127'b0000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000048000000000000000000000) 
14'h13f6 : LOC =         127'b0000000000000000000000000000000000010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000088000000000000000000000) 
14'h0369 : LOC =         127'b0000000000000000000000000000000000100001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000108000000000000000000000) 
14'h2257 : LOC =         127'b0000000000000000000000000000000001000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000208000000000000000000000) 
14'h235c : LOC =         127'b0000000000000000000000000000000010000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000408000000000000000000000) 
14'h214a : LOC =         127'b0000000000000000000000000000000100000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000808000000000000000000000) 
14'h2566 : LOC =         127'b0000000000000000000000000000001000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000001008000000000000000000000) 
14'h2d3e : LOC =         127'b0000000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000002008000000000000000000000) 
14'h3d8e : LOC =         127'b0000000000000000000000000000100000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000004008000000000000000000000) 
14'h1cee : LOC =         127'b0000000000000000000000000001000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000008008000000000000000000000) 
14'h1d59 : LOC =         127'b0000000000000000000000000010000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000010008000000000000000000000) 
14'h1e37 : LOC =         127'b0000000000000000000000000100000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000020008000000000000000000000) 
14'h18eb : LOC =         127'b0000000000000000000000001000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000040008000000000000000000000) 
14'h1553 : LOC =         127'b0000000000000000000000010000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000080008000000000000000000000) 
14'h0e23 : LOC =         127'b0000000000000000000000100000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000100008000000000000000000000) 
14'h38c3 : LOC =         127'b0000000000000000000001000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000200008000000000000000000000) 
14'h1674 : LOC =         127'b0000000000000000000010000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000400008000000000000000000000) 
14'h086d : LOC =         127'b0000000000000000000100000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000800008000000000000000000000) 
14'h345f : LOC =         127'b0000000000000000001000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00001000008000000000000000000000) 
14'h0f4c : LOC =         127'b0000000000000000010000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00002000008000000000000000000000) 
14'h3a1d : LOC =         127'b0000000000000000100000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00004000008000000000000000000000) 
14'h13c8 : LOC =         127'b0000000000000001000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00008000008000000000000000000000) 
14'h0315 : LOC =         127'b0000000000000010000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00010000008000000000000000000000) 
14'h22af : LOC =         127'b0000000000000100000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00020000008000000000000000000000) 
14'h22ac : LOC =         127'b0000000000001000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00040000008000000000000000000000) 
14'h22aa : LOC =         127'b0000000000010000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00080000008000000000000000000000) 
14'h22a6 : LOC =         127'b0000000000100000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00100000008000000000000000000000) 
14'h22be : LOC =         127'b0000000001000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00200000008000000000000000000000) 
14'h228e : LOC =         127'b0000000010000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00400000008000000000000000000000) 
14'h22ee : LOC =         127'b0000000100000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00800000008000000000000000000000) 
14'h222e : LOC =         127'b0000001000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x01000000008000000000000000000000) 
14'h23ae : LOC =         127'b0000010000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x02000000008000000000000000000000) 
14'h20ae : LOC =         127'b0000100000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x04000000008000000000000000000000) 
14'h26ae : LOC =         127'b0001000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x08000000008000000000000000000000) 
14'h2aae : LOC =         127'b0010000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x10000000008000000000000000000000) 
14'h32ae : LOC =         127'b0100000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x20000000008000000000000000000000) 
14'h02ae : LOC =         127'b1000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x40000000008000000000000000000000) 
14'h062b : LOC =         127'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // S (0x00000000010000000000000000000000) 
14'h0a7d : LOC =         127'b0000000000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000030000000000000000000000) 
14'h1e87 : LOC =         127'b0000000000000000000000000000000000001010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000050000000000000000000000) 
14'h3773 : LOC =         127'b0000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000090000000000000000000000) 
14'h27ec : LOC =         127'b0000000000000000000000000000000000100010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000110000000000000000000000) 
14'h06d2 : LOC =         127'b0000000000000000000000000000000001000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000210000000000000000000000) 
14'h07d9 : LOC =         127'b0000000000000000000000000000000010000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000410000000000000000000000) 
14'h05cf : LOC =         127'b0000000000000000000000000000000100000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000810000000000000000000000) 
14'h01e3 : LOC =         127'b0000000000000000000000000000001000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000001010000000000000000000000) 
14'h09bb : LOC =         127'b0000000000000000000000000000010000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000002010000000000000000000000) 
14'h190b : LOC =         127'b0000000000000000000000000000100000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000004010000000000000000000000) 
14'h386b : LOC =         127'b0000000000000000000000000001000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000008010000000000000000000000) 
14'h39dc : LOC =         127'b0000000000000000000000000010000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000010010000000000000000000000) 
14'h3ab2 : LOC =         127'b0000000000000000000000000100000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000020010000000000000000000000) 
14'h3c6e : LOC =         127'b0000000000000000000000001000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000040010000000000000000000000) 
14'h31d6 : LOC =         127'b0000000000000000000000010000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000080010000000000000000000000) 
14'h2aa6 : LOC =         127'b0000000000000000000000100000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000100010000000000000000000000) 
14'h1c46 : LOC =         127'b0000000000000000000001000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000200010000000000000000000000) 
14'h32f1 : LOC =         127'b0000000000000000000010000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000400010000000000000000000000) 
14'h2ce8 : LOC =         127'b0000000000000000000100000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000800010000000000000000000000) 
14'h10da : LOC =         127'b0000000000000000001000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00001000010000000000000000000000) 
14'h2bc9 : LOC =         127'b0000000000000000010000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00002000010000000000000000000000) 
14'h1e98 : LOC =         127'b0000000000000000100000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00004000010000000000000000000000) 
14'h374d : LOC =         127'b0000000000000001000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00008000010000000000000000000000) 
14'h2790 : LOC =         127'b0000000000000010000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00010000010000000000000000000000) 
14'h062a : LOC =         127'b0000000000000100000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00020000010000000000000000000000) 
14'h0629 : LOC =         127'b0000000000001000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00040000010000000000000000000000) 
14'h062f : LOC =         127'b0000000000010000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00080000010000000000000000000000) 
14'h0623 : LOC =         127'b0000000000100000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00100000010000000000000000000000) 
14'h063b : LOC =         127'b0000000001000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00200000010000000000000000000000) 
14'h060b : LOC =         127'b0000000010000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00400000010000000000000000000000) 
14'h066b : LOC =         127'b0000000100000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00800000010000000000000000000000) 
14'h06ab : LOC =         127'b0000001000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x01000000010000000000000000000000) 
14'h072b : LOC =         127'b0000010000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x02000000010000000000000000000000) 
14'h042b : LOC =         127'b0000100000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x04000000010000000000000000000000) 
14'h022b : LOC =         127'b0001000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x08000000010000000000000000000000) 
14'h0e2b : LOC =         127'b0010000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x10000000010000000000000000000000) 
14'h162b : LOC =         127'b0100000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x20000000010000000000000000000000) 
14'h262b : LOC =         127'b1000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x40000000010000000000000000000000) 
14'h0c56 : LOC =         127'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // S (0x00000000020000000000000000000000) 
14'h14fa : LOC =         127'b0000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000060000000000000000000000) 
14'h3d0e : LOC =         127'b0000000000000000000000000000000000010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x000000000a0000000000000000000000) 
14'h2d91 : LOC =         127'b0000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000120000000000000000000000) 
14'h0caf : LOC =         127'b0000000000000000000000000000000001000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000220000000000000000000000) 
14'h0da4 : LOC =         127'b0000000000000000000000000000000010000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000420000000000000000000000) 
14'h0fb2 : LOC =         127'b0000000000000000000000000000000100000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000820000000000000000000000) 
14'h0b9e : LOC =         127'b0000000000000000000000000000001000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000001020000000000000000000000) 
14'h03c6 : LOC =         127'b0000000000000000000000000000010000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000002020000000000000000000000) 
14'h1376 : LOC =         127'b0000000000000000000000000000100000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000004020000000000000000000000) 
14'h3216 : LOC =         127'b0000000000000000000000000001000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000008020000000000000000000000) 
14'h33a1 : LOC =         127'b0000000000000000000000000010000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000010020000000000000000000000) 
14'h30cf : LOC =         127'b0000000000000000000000000100000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000020020000000000000000000000) 
14'h3613 : LOC =         127'b0000000000000000000000001000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000040020000000000000000000000) 
14'h3bab : LOC =         127'b0000000000000000000000010000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000080020000000000000000000000) 
14'h20db : LOC =         127'b0000000000000000000000100000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000100020000000000000000000000) 
14'h163b : LOC =         127'b0000000000000000000001000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000200020000000000000000000000) 
14'h388c : LOC =         127'b0000000000000000000010000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000400020000000000000000000000) 
14'h2695 : LOC =         127'b0000000000000000000100000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000800020000000000000000000000) 
14'h1aa7 : LOC =         127'b0000000000000000001000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00001000020000000000000000000000) 
14'h21b4 : LOC =         127'b0000000000000000010000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00002000020000000000000000000000) 
14'h14e5 : LOC =         127'b0000000000000000100000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00004000020000000000000000000000) 
14'h3d30 : LOC =         127'b0000000000000001000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00008000020000000000000000000000) 
14'h2ded : LOC =         127'b0000000000000010000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00010000020000000000000000000000) 
14'h0c57 : LOC =         127'b0000000000000100000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00020000020000000000000000000000) 
14'h0c54 : LOC =         127'b0000000000001000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00040000020000000000000000000000) 
14'h0c52 : LOC =         127'b0000000000010000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00080000020000000000000000000000) 
14'h0c5e : LOC =         127'b0000000000100000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00100000020000000000000000000000) 
14'h0c46 : LOC =         127'b0000000001000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00200000020000000000000000000000) 
14'h0c76 : LOC =         127'b0000000010000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00400000020000000000000000000000) 
14'h0c16 : LOC =         127'b0000000100000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00800000020000000000000000000000) 
14'h0cd6 : LOC =         127'b0000001000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x01000000020000000000000000000000) 
14'h0d56 : LOC =         127'b0000010000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x02000000020000000000000000000000) 
14'h0e56 : LOC =         127'b0000100000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x04000000020000000000000000000000) 
14'h0856 : LOC =         127'b0001000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x08000000020000000000000000000000) 
14'h0456 : LOC =         127'b0010000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x10000000020000000000000000000000) 
14'h1c56 : LOC =         127'b0100000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x20000000020000000000000000000000) 
14'h2c56 : LOC =         127'b1000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x40000000020000000000000000000000) 
14'h18ac : LOC =         127'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // S (0x00000000040000000000000000000000) 
14'h29f4 : LOC =         127'b0000000000000000000000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x000000000c0000000000000000000000) 
14'h396b : LOC =         127'b0000000000000000000000000000000000101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000140000000000000000000000) 
14'h1855 : LOC =         127'b0000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000240000000000000000000000) 
14'h195e : LOC =         127'b0000000000000000000000000000000010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000440000000000000000000000) 
14'h1b48 : LOC =         127'b0000000000000000000000000000000100001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000840000000000000000000000) 
14'h1f64 : LOC =         127'b0000000000000000000000000000001000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000001040000000000000000000000) 
14'h173c : LOC =         127'b0000000000000000000000000000010000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000002040000000000000000000000) 
14'h078c : LOC =         127'b0000000000000000000000000000100000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000004040000000000000000000000) 
14'h26ec : LOC =         127'b0000000000000000000000000001000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000008040000000000000000000000) 
14'h275b : LOC =         127'b0000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000010040000000000000000000000) 
14'h2435 : LOC =         127'b0000000000000000000000000100000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000020040000000000000000000000) 
14'h22e9 : LOC =         127'b0000000000000000000000001000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000040040000000000000000000000) 
14'h2f51 : LOC =         127'b0000000000000000000000010000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000080040000000000000000000000) 
14'h3421 : LOC =         127'b0000000000000000000000100000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000100040000000000000000000000) 
14'h02c1 : LOC =         127'b0000000000000000000001000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000200040000000000000000000000) 
14'h2c76 : LOC =         127'b0000000000000000000010000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000400040000000000000000000000) 
14'h326f : LOC =         127'b0000000000000000000100000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000800040000000000000000000000) 
14'h0e5d : LOC =         127'b0000000000000000001000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00001000040000000000000000000000) 
14'h354e : LOC =         127'b0000000000000000010000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00002000040000000000000000000000) 
14'h001f : LOC =         127'b0000000000000000100000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00004000040000000000000000000000) 
14'h29ca : LOC =         127'b0000000000000001000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00008000040000000000000000000000) 
14'h3917 : LOC =         127'b0000000000000010000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00010000040000000000000000000000) 
14'h18ad : LOC =         127'b0000000000000100000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00020000040000000000000000000000) 
14'h18ae : LOC =         127'b0000000000001000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00040000040000000000000000000000) 
14'h18a8 : LOC =         127'b0000000000010000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00080000040000000000000000000000) 
14'h18a4 : LOC =         127'b0000000000100000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00100000040000000000000000000000) 
14'h18bc : LOC =         127'b0000000001000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00200000040000000000000000000000) 
14'h188c : LOC =         127'b0000000010000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00400000040000000000000000000000) 
14'h18ec : LOC =         127'b0000000100000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00800000040000000000000000000000) 
14'h182c : LOC =         127'b0000001000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x01000000040000000000000000000000) 
14'h19ac : LOC =         127'b0000010000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x02000000040000000000000000000000) 
14'h1aac : LOC =         127'b0000100000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x04000000040000000000000000000000) 
14'h1cac : LOC =         127'b0001000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x08000000040000000000000000000000) 
14'h10ac : LOC =         127'b0010000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x10000000040000000000000000000000) 
14'h08ac : LOC =         127'b0100000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x20000000040000000000000000000000) 
14'h38ac : LOC =         127'b1000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x40000000040000000000000000000000) 
14'h3158 : LOC =         127'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // S (0x00000000080000000000000000000000) 
14'h109f : LOC =         127'b0000000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000180000000000000000000000) 
14'h31a1 : LOC =         127'b0000000000000000000000000000000001010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000280000000000000000000000) 
14'h30aa : LOC =         127'b0000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000480000000000000000000000) 
14'h32bc : LOC =         127'b0000000000000000000000000000000100010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000880000000000000000000000) 
14'h3690 : LOC =         127'b0000000000000000000000000000001000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000001080000000000000000000000) 
14'h3ec8 : LOC =         127'b0000000000000000000000000000010000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000002080000000000000000000000) 
14'h2e78 : LOC =         127'b0000000000000000000000000000100000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000004080000000000000000000000) 
14'h0f18 : LOC =         127'b0000000000000000000000000001000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000008080000000000000000000000) 
14'h0eaf : LOC =         127'b0000000000000000000000000010000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000010080000000000000000000000) 
14'h0dc1 : LOC =         127'b0000000000000000000000000100000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000020080000000000000000000000) 
14'h0b1d : LOC =         127'b0000000000000000000000001000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000040080000000000000000000000) 
14'h06a5 : LOC =         127'b0000000000000000000000010000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000080080000000000000000000000) 
14'h1dd5 : LOC =         127'b0000000000000000000000100000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000100080000000000000000000000) 
14'h2b35 : LOC =         127'b0000000000000000000001000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000200080000000000000000000000) 
14'h0582 : LOC =         127'b0000000000000000000010000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000400080000000000000000000000) 
14'h1b9b : LOC =         127'b0000000000000000000100000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000800080000000000000000000000) 
14'h27a9 : LOC =         127'b0000000000000000001000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00001000080000000000000000000000) 
14'h1cba : LOC =         127'b0000000000000000010000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00002000080000000000000000000000) 
14'h29eb : LOC =         127'b0000000000000000100000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00004000080000000000000000000000) 
14'h003e : LOC =         127'b0000000000000001000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00008000080000000000000000000000) 
14'h10e3 : LOC =         127'b0000000000000010000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00010000080000000000000000000000) 
14'h3159 : LOC =         127'b0000000000000100000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00020000080000000000000000000000) 
14'h315a : LOC =         127'b0000000000001000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00040000080000000000000000000000) 
14'h315c : LOC =         127'b0000000000010000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00080000080000000000000000000000) 
14'h3150 : LOC =         127'b0000000000100000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00100000080000000000000000000000) 
14'h3148 : LOC =         127'b0000000001000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00200000080000000000000000000000) 
14'h3178 : LOC =         127'b0000000010000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00400000080000000000000000000000) 
14'h3118 : LOC =         127'b0000000100000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00800000080000000000000000000000) 
14'h31d8 : LOC =         127'b0000001000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x01000000080000000000000000000000) 
14'h3058 : LOC =         127'b0000010000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x02000000080000000000000000000000) 
14'h3358 : LOC =         127'b0000100000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x04000000080000000000000000000000) 
14'h3558 : LOC =         127'b0001000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x08000000080000000000000000000000) 
14'h3958 : LOC =         127'b0010000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x10000000080000000000000000000000) 
14'h2158 : LOC =         127'b0100000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x20000000080000000000000000000000) 
14'h1158 : LOC =         127'b1000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x40000000080000000000000000000000) 
14'h21c7 : LOC =         127'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // S (0x00000000100000000000000000000000) 
14'h213e : LOC =         127'b0000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000300000000000000000000000) 
14'h2035 : LOC =         127'b0000000000000000000000000000000010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000500000000000000000000000) 
14'h2223 : LOC =         127'b0000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000900000000000000000000000) 
14'h260f : LOC =         127'b0000000000000000000000000000001000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000001100000000000000000000000) 
14'h2e57 : LOC =         127'b0000000000000000000000000000010000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000002100000000000000000000000) 
14'h3ee7 : LOC =         127'b0000000000000000000000000000100000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000004100000000000000000000000) 
14'h1f87 : LOC =         127'b0000000000000000000000000001000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000008100000000000000000000000) 
14'h1e30 : LOC =         127'b0000000000000000000000000010000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000010100000000000000000000000) 
14'h1d5e : LOC =         127'b0000000000000000000000000100000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000020100000000000000000000000) 
14'h1b82 : LOC =         127'b0000000000000000000000001000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000040100000000000000000000000) 
14'h163a : LOC =         127'b0000000000000000000000010000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000080100000000000000000000000) 
14'h0d4a : LOC =         127'b0000000000000000000000100000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000100100000000000000000000000) 
14'h3baa : LOC =         127'b0000000000000000000001000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000200100000000000000000000000) 
14'h151d : LOC =         127'b0000000000000000000010000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000400100000000000000000000000) 
14'h0b04 : LOC =         127'b0000000000000000000100000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000800100000000000000000000000) 
14'h3736 : LOC =         127'b0000000000000000001000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00001000100000000000000000000000) 
14'h0c25 : LOC =         127'b0000000000000000010000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00002000100000000000000000000000) 
14'h3974 : LOC =         127'b0000000000000000100000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00004000100000000000000000000000) 
14'h10a1 : LOC =         127'b0000000000000001000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00008000100000000000000000000000) 
14'h007c : LOC =         127'b0000000000000010000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00010000100000000000000000000000) 
14'h21c6 : LOC =         127'b0000000000000100000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00020000100000000000000000000000) 
14'h21c5 : LOC =         127'b0000000000001000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00040000100000000000000000000000) 
14'h21c3 : LOC =         127'b0000000000010000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00080000100000000000000000000000) 
14'h21cf : LOC =         127'b0000000000100000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00100000100000000000000000000000) 
14'h21d7 : LOC =         127'b0000000001000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00200000100000000000000000000000) 
14'h21e7 : LOC =         127'b0000000010000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00400000100000000000000000000000) 
14'h2187 : LOC =         127'b0000000100000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00800000100000000000000000000000) 
14'h2147 : LOC =         127'b0000001000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x01000000100000000000000000000000) 
14'h20c7 : LOC =         127'b0000010000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x02000000100000000000000000000000) 
14'h23c7 : LOC =         127'b0000100000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x04000000100000000000000000000000) 
14'h25c7 : LOC =         127'b0001000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x08000000100000000000000000000000) 
14'h29c7 : LOC =         127'b0010000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x10000000100000000000000000000000) 
14'h31c7 : LOC =         127'b0100000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x20000000100000000000000000000000) 
14'h01c7 : LOC =         127'b1000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x40000000100000000000000000000000) 
14'h00f9 : LOC =         127'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // S (0x00000000200000000000000000000000) 
14'h010b : LOC =         127'b0000000000000000000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000600000000000000000000000) 
14'h031d : LOC =         127'b0000000000000000000000000000000101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000a00000000000000000000000) 
14'h0731 : LOC =         127'b0000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000001200000000000000000000000) 
14'h0f69 : LOC =         127'b0000000000000000000000000000010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000002200000000000000000000000) 
14'h1fd9 : LOC =         127'b0000000000000000000000000000100001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000004200000000000000000000000) 
14'h3eb9 : LOC =         127'b0000000000000000000000000001000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000008200000000000000000000000) 
14'h3f0e : LOC =         127'b0000000000000000000000000010000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000010200000000000000000000000) 
14'h3c60 : LOC =         127'b0000000000000000000000000100000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000020200000000000000000000000) 
14'h3abc : LOC =         127'b0000000000000000000000001000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000040200000000000000000000000) 
14'h3704 : LOC =         127'b0000000000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000080200000000000000000000000) 
14'h2c74 : LOC =         127'b0000000000000000000000100000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000100200000000000000000000000) 
14'h1a94 : LOC =         127'b0000000000000000000001000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000200200000000000000000000000) 
14'h3423 : LOC =         127'b0000000000000000000010000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000400200000000000000000000000) 
14'h2a3a : LOC =         127'b0000000000000000000100000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000800200000000000000000000000) 
14'h1608 : LOC =         127'b0000000000000000001000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00001000200000000000000000000000) 
14'h2d1b : LOC =         127'b0000000000000000010000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00002000200000000000000000000000) 
14'h184a : LOC =         127'b0000000000000000100000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00004000200000000000000000000000) 
14'h319f : LOC =         127'b0000000000000001000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00008000200000000000000000000000) 
14'h2142 : LOC =         127'b0000000000000010000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00010000200000000000000000000000) 
14'h00f8 : LOC =         127'b0000000000000100000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00020000200000000000000000000000) 
14'h00fb : LOC =         127'b0000000000001000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00040000200000000000000000000000) 
14'h00fd : LOC =         127'b0000000000010000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00080000200000000000000000000000) 
14'h00f1 : LOC =         127'b0000000000100000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00100000200000000000000000000000) 
14'h00e9 : LOC =         127'b0000000001000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00200000200000000000000000000000) 
14'h00d9 : LOC =         127'b0000000010000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00400000200000000000000000000000) 
14'h00b9 : LOC =         127'b0000000100000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00800000200000000000000000000000) 
14'h0079 : LOC =         127'b0000001000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x01000000200000000000000000000000) 
14'h01f9 : LOC =         127'b0000010000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x02000000200000000000000000000000) 
14'h02f9 : LOC =         127'b0000100000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x04000000200000000000000000000000) 
14'h04f9 : LOC =         127'b0001000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x08000000200000000000000000000000) 
14'h08f9 : LOC =         127'b0010000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x10000000200000000000000000000000) 
14'h10f9 : LOC =         127'b0100000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x20000000200000000000000000000000) 
14'h20f9 : LOC =         127'b1000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x40000000200000000000000000000000) 
14'h01f2 : LOC =         127'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // S (0x00000000400000000000000000000000) 
14'h0216 : LOC =         127'b0000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000000c00000000000000000000000) 
14'h063a : LOC =         127'b0000000000000000000000000000001010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000001400000000000000000000000) 
14'h0e62 : LOC =         127'b0000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000002400000000000000000000000) 
14'h1ed2 : LOC =         127'b0000000000000000000000000000100010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000004400000000000000000000000) 
14'h3fb2 : LOC =         127'b0000000000000000000000000001000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000008400000000000000000000000) 
14'h3e05 : LOC =         127'b0000000000000000000000000010000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000010400000000000000000000000) 
14'h3d6b : LOC =         127'b0000000000000000000000000100000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000020400000000000000000000000) 
14'h3bb7 : LOC =         127'b0000000000000000000000001000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000040400000000000000000000000) 
14'h360f : LOC =         127'b0000000000000000000000010000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000080400000000000000000000000) 
14'h2d7f : LOC =         127'b0000000000000000000000100000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000100400000000000000000000000) 
14'h1b9f : LOC =         127'b0000000000000000000001000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000200400000000000000000000000) 
14'h3528 : LOC =         127'b0000000000000000000010000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000400400000000000000000000000) 
14'h2b31 : LOC =         127'b0000000000000000000100000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000800400000000000000000000000) 
14'h1703 : LOC =         127'b0000000000000000001000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00001000400000000000000000000000) 
14'h2c10 : LOC =         127'b0000000000000000010000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00002000400000000000000000000000) 
14'h1941 : LOC =         127'b0000000000000000100000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00004000400000000000000000000000) 
14'h3094 : LOC =         127'b0000000000000001000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00008000400000000000000000000000) 
14'h2049 : LOC =         127'b0000000000000010000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00010000400000000000000000000000) 
14'h01f3 : LOC =         127'b0000000000000100000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00020000400000000000000000000000) 
14'h01f0 : LOC =         127'b0000000000001000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00040000400000000000000000000000) 
14'h01f6 : LOC =         127'b0000000000010000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00080000400000000000000000000000) 
14'h01fa : LOC =         127'b0000000000100000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00100000400000000000000000000000) 
14'h01e2 : LOC =         127'b0000000001000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00200000400000000000000000000000) 
14'h01d2 : LOC =         127'b0000000010000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00400000400000000000000000000000) 
14'h01b2 : LOC =         127'b0000000100000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00800000400000000000000000000000) 
14'h0172 : LOC =         127'b0000001000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x01000000400000000000000000000000) 
14'h00f2 : LOC =         127'b0000010000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x02000000400000000000000000000000) 
14'h03f2 : LOC =         127'b0000100000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x04000000400000000000000000000000) 
14'h05f2 : LOC =         127'b0001000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x08000000400000000000000000000000) 
14'h09f2 : LOC =         127'b0010000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x10000000400000000000000000000000) 
14'h11f2 : LOC =         127'b0100000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x20000000400000000000000000000000) 
14'h21f2 : LOC =         127'b1000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x40000000400000000000000000000000) 
14'h03e4 : LOC =         127'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // S (0x00000000800000000000000000000000) 
14'h042c : LOC =         127'b0000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000001800000000000000000000000) 
14'h0c74 : LOC =         127'b0000000000000000000000000000010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000002800000000000000000000000) 
14'h1cc4 : LOC =         127'b0000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000004800000000000000000000000) 
14'h3da4 : LOC =         127'b0000000000000000000000000001000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000008800000000000000000000000) 
14'h3c13 : LOC =         127'b0000000000000000000000000010000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000010800000000000000000000000) 
14'h3f7d : LOC =         127'b0000000000000000000000000100000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000020800000000000000000000000) 
14'h39a1 : LOC =         127'b0000000000000000000000001000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000040800000000000000000000000) 
14'h3419 : LOC =         127'b0000000000000000000000010000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000080800000000000000000000000) 
14'h2f69 : LOC =         127'b0000000000000000000000100000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000100800000000000000000000000) 
14'h1989 : LOC =         127'b0000000000000000000001000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000200800000000000000000000000) 
14'h373e : LOC =         127'b0000000000000000000010000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000400800000000000000000000000) 
14'h2927 : LOC =         127'b0000000000000000000100000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000800800000000000000000000000) 
14'h1515 : LOC =         127'b0000000000000000001000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00001000800000000000000000000000) 
14'h2e06 : LOC =         127'b0000000000000000010000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00002000800000000000000000000000) 
14'h1b57 : LOC =         127'b0000000000000000100000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00004000800000000000000000000000) 
14'h3282 : LOC =         127'b0000000000000001000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00008000800000000000000000000000) 
14'h225f : LOC =         127'b0000000000000010000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00010000800000000000000000000000) 
14'h03e5 : LOC =         127'b0000000000000100000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00020000800000000000000000000000) 
14'h03e6 : LOC =         127'b0000000000001000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00040000800000000000000000000000) 
14'h03e0 : LOC =         127'b0000000000010000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00080000800000000000000000000000) 
14'h03ec : LOC =         127'b0000000000100000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00100000800000000000000000000000) 
14'h03f4 : LOC =         127'b0000000001000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00200000800000000000000000000000) 
14'h03c4 : LOC =         127'b0000000010000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00400000800000000000000000000000) 
14'h03a4 : LOC =         127'b0000000100000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00800000800000000000000000000000) 
14'h0364 : LOC =         127'b0000001000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x01000000800000000000000000000000) 
14'h02e4 : LOC =         127'b0000010000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x02000000800000000000000000000000) 
14'h01e4 : LOC =         127'b0000100000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x04000000800000000000000000000000) 
14'h07e4 : LOC =         127'b0001000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x08000000800000000000000000000000) 
14'h0be4 : LOC =         127'b0010000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x10000000800000000000000000000000) 
14'h13e4 : LOC =         127'b0100000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x20000000800000000000000000000000) 
14'h23e4 : LOC =         127'b1000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x40000000800000000000000000000000) 
14'h07c8 : LOC =         127'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // S (0x00000001000000000000000000000000) 
14'h0858 : LOC =         127'b0000000000000000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000003000000000000000000000000) 
14'h18e8 : LOC =         127'b0000000000000000000000000000101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000005000000000000000000000000) 
14'h3988 : LOC =         127'b0000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000009000000000000000000000000) 
14'h383f : LOC =         127'b0000000000000000000000000010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000011000000000000000000000000) 
14'h3b51 : LOC =         127'b0000000000000000000000000100001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000021000000000000000000000000) 
14'h3d8d : LOC =         127'b0000000000000000000000001000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000041000000000000000000000000) 
14'h3035 : LOC =         127'b0000000000000000000000010000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000081000000000000000000000000) 
14'h2b45 : LOC =         127'b0000000000000000000000100000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000101000000000000000000000000) 
14'h1da5 : LOC =         127'b0000000000000000000001000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000201000000000000000000000000) 
14'h3312 : LOC =         127'b0000000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000401000000000000000000000000) 
14'h2d0b : LOC =         127'b0000000000000000000100000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000801000000000000000000000000) 
14'h1139 : LOC =         127'b0000000000000000001000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00001001000000000000000000000000) 
14'h2a2a : LOC =         127'b0000000000000000010000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00002001000000000000000000000000) 
14'h1f7b : LOC =         127'b0000000000000000100000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00004001000000000000000000000000) 
14'h36ae : LOC =         127'b0000000000000001000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00008001000000000000000000000000) 
14'h2673 : LOC =         127'b0000000000000010000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00010001000000000000000000000000) 
14'h07c9 : LOC =         127'b0000000000000100000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00020001000000000000000000000000) 
14'h07ca : LOC =         127'b0000000000001000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00040001000000000000000000000000) 
14'h07cc : LOC =         127'b0000000000010000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00080001000000000000000000000000) 
14'h07c0 : LOC =         127'b0000000000100000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00100001000000000000000000000000) 
14'h07d8 : LOC =         127'b0000000001000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00200001000000000000000000000000) 
14'h07e8 : LOC =         127'b0000000010000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00400001000000000000000000000000) 
14'h0788 : LOC =         127'b0000000100000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00800001000000000000000000000000) 
14'h0748 : LOC =         127'b0000001000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x01000001000000000000000000000000) 
14'h06c8 : LOC =         127'b0000010000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x02000001000000000000000000000000) 
14'h05c8 : LOC =         127'b0000100000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x04000001000000000000000000000000) 
14'h03c8 : LOC =         127'b0001000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x08000001000000000000000000000000) 
14'h0fc8 : LOC =         127'b0010000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x10000001000000000000000000000000) 
14'h17c8 : LOC =         127'b0100000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x20000001000000000000000000000000) 
14'h27c8 : LOC =         127'b1000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x40000001000000000000000000000000) 
14'h0f90 : LOC =         127'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // S (0x00000002000000000000000000000000) 
14'h10b0 : LOC =         127'b0000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000006000000000000000000000000) 
14'h31d0 : LOC =         127'b0000000000000000000000000001010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x0000000a000000000000000000000000) 
14'h3067 : LOC =         127'b0000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000012000000000000000000000000) 
14'h3309 : LOC =         127'b0000000000000000000000000100010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000022000000000000000000000000) 
14'h35d5 : LOC =         127'b0000000000000000000000001000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000042000000000000000000000000) 
14'h386d : LOC =         127'b0000000000000000000000010000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000082000000000000000000000000) 
14'h231d : LOC =         127'b0000000000000000000000100000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000102000000000000000000000000) 
14'h15fd : LOC =         127'b0000000000000000000001000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000202000000000000000000000000) 
14'h3b4a : LOC =         127'b0000000000000000000010000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000402000000000000000000000000) 
14'h2553 : LOC =         127'b0000000000000000000100000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000802000000000000000000000000) 
14'h1961 : LOC =         127'b0000000000000000001000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00001002000000000000000000000000) 
14'h2272 : LOC =         127'b0000000000000000010000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00002002000000000000000000000000) 
14'h1723 : LOC =         127'b0000000000000000100000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00004002000000000000000000000000) 
14'h3ef6 : LOC =         127'b0000000000000001000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00008002000000000000000000000000) 
14'h2e2b : LOC =         127'b0000000000000010000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00010002000000000000000000000000) 
14'h0f91 : LOC =         127'b0000000000000100000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00020002000000000000000000000000) 
14'h0f92 : LOC =         127'b0000000000001000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00040002000000000000000000000000) 
14'h0f94 : LOC =         127'b0000000000010000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00080002000000000000000000000000) 
14'h0f98 : LOC =         127'b0000000000100000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00100002000000000000000000000000) 
14'h0f80 : LOC =         127'b0000000001000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00200002000000000000000000000000) 
14'h0fb0 : LOC =         127'b0000000010000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00400002000000000000000000000000) 
14'h0fd0 : LOC =         127'b0000000100000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00800002000000000000000000000000) 
14'h0f10 : LOC =         127'b0000001000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x01000002000000000000000000000000) 
14'h0e90 : LOC =         127'b0000010000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x02000002000000000000000000000000) 
14'h0d90 : LOC =         127'b0000100000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x04000002000000000000000000000000) 
14'h0b90 : LOC =         127'b0001000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x08000002000000000000000000000000) 
14'h0790 : LOC =         127'b0010000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x10000002000000000000000000000000) 
14'h1f90 : LOC =         127'b0100000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x20000002000000000000000000000000) 
14'h2f90 : LOC =         127'b1000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x40000002000000000000000000000000) 
14'h1f20 : LOC =         127'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // S (0x00000004000000000000000000000000) 
14'h2160 : LOC =         127'b0000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x0000000c000000000000000000000000) 
14'h20d7 : LOC =         127'b0000000000000000000000000010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000014000000000000000000000000) 
14'h23b9 : LOC =         127'b0000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000024000000000000000000000000) 
14'h2565 : LOC =         127'b0000000000000000000000001000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000044000000000000000000000000) 
14'h28dd : LOC =         127'b0000000000000000000000010000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000084000000000000000000000000) 
14'h33ad : LOC =         127'b0000000000000000000000100000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000104000000000000000000000000) 
14'h054d : LOC =         127'b0000000000000000000001000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000204000000000000000000000000) 
14'h2bfa : LOC =         127'b0000000000000000000010000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000404000000000000000000000000) 
14'h35e3 : LOC =         127'b0000000000000000000100000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000804000000000000000000000000) 
14'h09d1 : LOC =         127'b0000000000000000001000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00001004000000000000000000000000) 
14'h32c2 : LOC =         127'b0000000000000000010000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00002004000000000000000000000000) 
14'h0793 : LOC =         127'b0000000000000000100000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00004004000000000000000000000000) 
14'h2e46 : LOC =         127'b0000000000000001000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00008004000000000000000000000000) 
14'h3e9b : LOC =         127'b0000000000000010000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00010004000000000000000000000000) 
14'h1f21 : LOC =         127'b0000000000000100000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00020004000000000000000000000000) 
14'h1f22 : LOC =         127'b0000000000001000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00040004000000000000000000000000) 
14'h1f24 : LOC =         127'b0000000000010000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00080004000000000000000000000000) 
14'h1f28 : LOC =         127'b0000000000100000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00100004000000000000000000000000) 
14'h1f30 : LOC =         127'b0000000001000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00200004000000000000000000000000) 
14'h1f00 : LOC =         127'b0000000010000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00400004000000000000000000000000) 
14'h1f60 : LOC =         127'b0000000100000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00800004000000000000000000000000) 
14'h1fa0 : LOC =         127'b0000001000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x01000004000000000000000000000000) 
14'h1e20 : LOC =         127'b0000010000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x02000004000000000000000000000000) 
14'h1d20 : LOC =         127'b0000100000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x04000004000000000000000000000000) 
14'h1b20 : LOC =         127'b0001000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x08000004000000000000000000000000) 
14'h1720 : LOC =         127'b0010000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x10000004000000000000000000000000) 
14'h0f20 : LOC =         127'b0100000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x20000004000000000000000000000000) 
14'h3f20 : LOC =         127'b1000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x40000004000000000000000000000000) 
14'h3e40 : LOC =         127'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // S (0x00000008000000000000000000000000) 
14'h01b7 : LOC =         127'b0000000000000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000018000000000000000000000000) 
14'h02d9 : LOC =         127'b0000000000000000000000000101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000028000000000000000000000000) 
14'h0405 : LOC =         127'b0000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000048000000000000000000000000) 
14'h09bd : LOC =         127'b0000000000000000000000010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000088000000000000000000000000) 
14'h12cd : LOC =         127'b0000000000000000000000100001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000108000000000000000000000000) 
14'h242d : LOC =         127'b0000000000000000000001000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000208000000000000000000000000) 
14'h0a9a : LOC =         127'b0000000000000000000010000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000408000000000000000000000000) 
14'h1483 : LOC =         127'b0000000000000000000100000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000808000000000000000000000000) 
14'h28b1 : LOC =         127'b0000000000000000001000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00001008000000000000000000000000) 
14'h13a2 : LOC =         127'b0000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00002008000000000000000000000000) 
14'h26f3 : LOC =         127'b0000000000000000100000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00004008000000000000000000000000) 
14'h0f26 : LOC =         127'b0000000000000001000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00008008000000000000000000000000) 
14'h1ffb : LOC =         127'b0000000000000010000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00010008000000000000000000000000) 
14'h3e41 : LOC =         127'b0000000000000100000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00020008000000000000000000000000) 
14'h3e42 : LOC =         127'b0000000000001000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00040008000000000000000000000000) 
14'h3e44 : LOC =         127'b0000000000010000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00080008000000000000000000000000) 
14'h3e48 : LOC =         127'b0000000000100000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00100008000000000000000000000000) 
14'h3e50 : LOC =         127'b0000000001000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00200008000000000000000000000000) 
14'h3e60 : LOC =         127'b0000000010000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00400008000000000000000000000000) 
14'h3e00 : LOC =         127'b0000000100000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00800008000000000000000000000000) 
14'h3ec0 : LOC =         127'b0000001000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x01000008000000000000000000000000) 
14'h3f40 : LOC =         127'b0000010000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x02000008000000000000000000000000) 
14'h3c40 : LOC =         127'b0000100000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x04000008000000000000000000000000) 
14'h3a40 : LOC =         127'b0001000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x08000008000000000000000000000000) 
14'h3640 : LOC =         127'b0010000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x10000008000000000000000000000000) 
14'h2e40 : LOC =         127'b0100000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x20000008000000000000000000000000) 
14'h1e40 : LOC =         127'b1000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x40000008000000000000000000000000) 
14'h3ff7 : LOC =         127'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // S (0x00000010000000000000000000000000) 
14'h036e : LOC =         127'b0000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000030000000000000000000000000) 
14'h05b2 : LOC =         127'b0000000000000000000000001010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000050000000000000000000000000) 
14'h080a : LOC =         127'b0000000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000090000000000000000000000000) 
14'h137a : LOC =         127'b0000000000000000000000100010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000110000000000000000000000000) 
14'h259a : LOC =         127'b0000000000000000000001000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000210000000000000000000000000) 
14'h0b2d : LOC =         127'b0000000000000000000010000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000410000000000000000000000000) 
14'h1534 : LOC =         127'b0000000000000000000100000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000810000000000000000000000000) 
14'h2906 : LOC =         127'b0000000000000000001000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00001010000000000000000000000000) 
14'h1215 : LOC =         127'b0000000000000000010000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00002010000000000000000000000000) 
14'h2744 : LOC =         127'b0000000000000000100000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00004010000000000000000000000000) 
14'h0e91 : LOC =         127'b0000000000000001000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00008010000000000000000000000000) 
14'h1e4c : LOC =         127'b0000000000000010000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00010010000000000000000000000000) 
14'h3ff6 : LOC =         127'b0000000000000100000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00020010000000000000000000000000) 
14'h3ff5 : LOC =         127'b0000000000001000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00040010000000000000000000000000) 
14'h3ff3 : LOC =         127'b0000000000010000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00080010000000000000000000000000) 
14'h3fff : LOC =         127'b0000000000100000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00100010000000000000000000000000) 
14'h3fe7 : LOC =         127'b0000000001000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00200010000000000000000000000000) 
14'h3fd7 : LOC =         127'b0000000010000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00400010000000000000000000000000) 
14'h3fb7 : LOC =         127'b0000000100000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00800010000000000000000000000000) 
14'h3f77 : LOC =         127'b0000001000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x01000010000000000000000000000000) 
14'h3ef7 : LOC =         127'b0000010000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x02000010000000000000000000000000) 
14'h3df7 : LOC =         127'b0000100000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x04000010000000000000000000000000) 
14'h3bf7 : LOC =         127'b0001000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x08000010000000000000000000000000) 
14'h37f7 : LOC =         127'b0010000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x10000010000000000000000000000000) 
14'h2ff7 : LOC =         127'b0100000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x20000010000000000000000000000000) 
14'h1ff7 : LOC =         127'b1000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x40000010000000000000000000000000) 
14'h3c99 : LOC =         127'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // S (0x00000020000000000000000000000000) 
14'h06dc : LOC =         127'b0000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000060000000000000000000000000) 
14'h0b64 : LOC =         127'b0000000000000000000000010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x000000a0000000000000000000000000) 
14'h1014 : LOC =         127'b0000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000120000000000000000000000000) 
14'h26f4 : LOC =         127'b0000000000000000000001000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000220000000000000000000000000) 
14'h0843 : LOC =         127'b0000000000000000000010000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000420000000000000000000000000) 
14'h165a : LOC =         127'b0000000000000000000100000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000820000000000000000000000000) 
14'h2a68 : LOC =         127'b0000000000000000001000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00001020000000000000000000000000) 
14'h117b : LOC =         127'b0000000000000000010000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00002020000000000000000000000000) 
14'h242a : LOC =         127'b0000000000000000100000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00004020000000000000000000000000) 
14'h0dff : LOC =         127'b0000000000000001000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00008020000000000000000000000000) 
14'h1d22 : LOC =         127'b0000000000000010000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00010020000000000000000000000000) 
14'h3c98 : LOC =         127'b0000000000000100000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00020020000000000000000000000000) 
14'h3c9b : LOC =         127'b0000000000001000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00040020000000000000000000000000) 
14'h3c9d : LOC =         127'b0000000000010000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00080020000000000000000000000000) 
14'h3c91 : LOC =         127'b0000000000100000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00100020000000000000000000000000) 
14'h3c89 : LOC =         127'b0000000001000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00200020000000000000000000000000) 
14'h3cb9 : LOC =         127'b0000000010000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00400020000000000000000000000000) 
14'h3cd9 : LOC =         127'b0000000100000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00800020000000000000000000000000) 
14'h3c19 : LOC =         127'b0000001000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x01000020000000000000000000000000) 
14'h3d99 : LOC =         127'b0000010000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x02000020000000000000000000000000) 
14'h3e99 : LOC =         127'b0000100000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x04000020000000000000000000000000) 
14'h3899 : LOC =         127'b0001000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x08000020000000000000000000000000) 
14'h3499 : LOC =         127'b0010000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x10000020000000000000000000000000) 
14'h2c99 : LOC =         127'b0100000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x20000020000000000000000000000000) 
14'h1c99 : LOC =         127'b1000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x40000020000000000000000000000000) 
14'h3a45 : LOC =         127'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // S (0x00000040000000000000000000000000) 
14'h0db8 : LOC =         127'b0000000000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x000000c0000000000000000000000000) 
14'h16c8 : LOC =         127'b0000000000000000000000101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000140000000000000000000000000) 
14'h2028 : LOC =         127'b0000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000240000000000000000000000000) 
14'h0e9f : LOC =         127'b0000000000000000000010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000440000000000000000000000000) 
14'h1086 : LOC =         127'b0000000000000000000100001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000840000000000000000000000000) 
14'h2cb4 : LOC =         127'b0000000000000000001000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00001040000000000000000000000000) 
14'h17a7 : LOC =         127'b0000000000000000010000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00002040000000000000000000000000) 
14'h22f6 : LOC =         127'b0000000000000000100000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00004040000000000000000000000000) 
14'h0b23 : LOC =         127'b0000000000000001000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00008040000000000000000000000000) 
14'h1bfe : LOC =         127'b0000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00010040000000000000000000000000) 
14'h3a44 : LOC =         127'b0000000000000100000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00020040000000000000000000000000) 
14'h3a47 : LOC =         127'b0000000000001000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00040040000000000000000000000000) 
14'h3a41 : LOC =         127'b0000000000010000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00080040000000000000000000000000) 
14'h3a4d : LOC =         127'b0000000000100000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00100040000000000000000000000000) 
14'h3a55 : LOC =         127'b0000000001000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00200040000000000000000000000000) 
14'h3a65 : LOC =         127'b0000000010000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00400040000000000000000000000000) 
14'h3a05 : LOC =         127'b0000000100000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00800040000000000000000000000000) 
14'h3ac5 : LOC =         127'b0000001000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x01000040000000000000000000000000) 
14'h3b45 : LOC =         127'b0000010000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x02000040000000000000000000000000) 
14'h3845 : LOC =         127'b0000100000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x04000040000000000000000000000000) 
14'h3e45 : LOC =         127'b0001000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x08000040000000000000000000000000) 
14'h3245 : LOC =         127'b0010000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x10000040000000000000000000000000) 
14'h2a45 : LOC =         127'b0100000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x20000040000000000000000000000000) 
14'h1a45 : LOC =         127'b1000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x40000040000000000000000000000000) 
14'h37fd : LOC =         127'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // S (0x00000080000000000000000000000000) 
14'h1b70 : LOC =         127'b0000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000180000000000000000000000000) 
14'h2d90 : LOC =         127'b0000000000000000000001010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000280000000000000000000000000) 
14'h0327 : LOC =         127'b0000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000480000000000000000000000000) 
14'h1d3e : LOC =         127'b0000000000000000000100010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000880000000000000000000000000) 
14'h210c : LOC =         127'b0000000000000000001000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00001080000000000000000000000000) 
14'h1a1f : LOC =         127'b0000000000000000010000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00002080000000000000000000000000) 
14'h2f4e : LOC =         127'b0000000000000000100000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00004080000000000000000000000000) 
14'h069b : LOC =         127'b0000000000000001000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00008080000000000000000000000000) 
14'h1646 : LOC =         127'b0000000000000010000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00010080000000000000000000000000) 
14'h37fc : LOC =         127'b0000000000000100000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00020080000000000000000000000000) 
14'h37ff : LOC =         127'b0000000000001000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00040080000000000000000000000000) 
14'h37f9 : LOC =         127'b0000000000010000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00080080000000000000000000000000) 
14'h37f5 : LOC =         127'b0000000000100000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00100080000000000000000000000000) 
14'h37ed : LOC =         127'b0000000001000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00200080000000000000000000000000) 
14'h37dd : LOC =         127'b0000000010000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00400080000000000000000000000000) 
14'h37bd : LOC =         127'b0000000100000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00800080000000000000000000000000) 
14'h377d : LOC =         127'b0000001000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x01000080000000000000000000000000) 
14'h36fd : LOC =         127'b0000010000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x02000080000000000000000000000000) 
14'h35fd : LOC =         127'b0000100000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x04000080000000000000000000000000) 
14'h33fd : LOC =         127'b0001000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x08000080000000000000000000000000) 
14'h3ffd : LOC =         127'b0010000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x10000080000000000000000000000000) 
14'h27fd : LOC =         127'b0100000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x20000080000000000000000000000000) 
14'h17fd : LOC =         127'b1000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x40000080000000000000000000000000) 
14'h2c8d : LOC =         127'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // S (0x00000100000000000000000000000000) 
14'h36e0 : LOC =         127'b0000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000300000000000000000000000000) 
14'h1857 : LOC =         127'b0000000000000000000010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000500000000000000000000000000) 
14'h064e : LOC =         127'b0000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000900000000000000000000000000) 
14'h3a7c : LOC =         127'b0000000000000000001000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00001100000000000000000000000000) 
14'h016f : LOC =         127'b0000000000000000010000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00002100000000000000000000000000) 
14'h343e : LOC =         127'b0000000000000000100000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00004100000000000000000000000000) 
14'h1deb : LOC =         127'b0000000000000001000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00008100000000000000000000000000) 
14'h0d36 : LOC =         127'b0000000000000010000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00010100000000000000000000000000) 
14'h2c8c : LOC =         127'b0000000000000100000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00020100000000000000000000000000) 
14'h2c8f : LOC =         127'b0000000000001000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00040100000000000000000000000000) 
14'h2c89 : LOC =         127'b0000000000010000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00080100000000000000000000000000) 
14'h2c85 : LOC =         127'b0000000000100000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00100100000000000000000000000000) 
14'h2c9d : LOC =         127'b0000000001000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00200100000000000000000000000000) 
14'h2cad : LOC =         127'b0000000010000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00400100000000000000000000000000) 
14'h2ccd : LOC =         127'b0000000100000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00800100000000000000000000000000) 
14'h2c0d : LOC =         127'b0000001000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x01000100000000000000000000000000) 
14'h2d8d : LOC =         127'b0000010000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x02000100000000000000000000000000) 
14'h2e8d : LOC =         127'b0000100000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x04000100000000000000000000000000) 
14'h288d : LOC =         127'b0001000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x08000100000000000000000000000000) 
14'h248d : LOC =         127'b0010000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x10000100000000000000000000000000) 
14'h3c8d : LOC =         127'b0100000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x20000100000000000000000000000000) 
14'h0c8d : LOC =         127'b1000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x40000100000000000000000000000000) 
14'h1a6d : LOC =         127'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // S (0x00000200000000000000000000000000) 
14'h2eb7 : LOC =         127'b0000000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000600000000000000000000000000) 
14'h30ae : LOC =         127'b0000000000000000000101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000a00000000000000000000000000) 
14'h0c9c : LOC =         127'b0000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00001200000000000000000000000000) 
14'h378f : LOC =         127'b0000000000000000010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00002200000000000000000000000000) 
14'h02de : LOC =         127'b0000000000000000100001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00004200000000000000000000000000) 
14'h2b0b : LOC =         127'b0000000000000001000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00008200000000000000000000000000) 
14'h3bd6 : LOC =         127'b0000000000000010000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00010200000000000000000000000000) 
14'h1a6c : LOC =         127'b0000000000000100000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00020200000000000000000000000000) 
14'h1a6f : LOC =         127'b0000000000001000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00040200000000000000000000000000) 
14'h1a69 : LOC =         127'b0000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00080200000000000000000000000000) 
14'h1a65 : LOC =         127'b0000000000100000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00100200000000000000000000000000) 
14'h1a7d : LOC =         127'b0000000001000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00200200000000000000000000000000) 
14'h1a4d : LOC =         127'b0000000010000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00400200000000000000000000000000) 
14'h1a2d : LOC =         127'b0000000100000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00800200000000000000000000000000) 
14'h1aed : LOC =         127'b0000001000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x01000200000000000000000000000000) 
14'h1b6d : LOC =         127'b0000010000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x02000200000000000000000000000000) 
14'h186d : LOC =         127'b0000100000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x04000200000000000000000000000000) 
14'h1e6d : LOC =         127'b0001000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x08000200000000000000000000000000) 
14'h126d : LOC =         127'b0010000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x10000200000000000000000000000000) 
14'h0a6d : LOC =         127'b0100000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x20000200000000000000000000000000) 
14'h3a6d : LOC =         127'b1000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x40000200000000000000000000000000) 
14'h34da : LOC =         127'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // S (0x00000400000000000000000000000000) 
14'h1e19 : LOC =         127'b0000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00000c00000000000000000000000000) 
14'h222b : LOC =         127'b0000000000000000001010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00001400000000000000000000000000) 
14'h1938 : LOC =         127'b0000000000000000010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00002400000000000000000000000000) 
14'h2c69 : LOC =         127'b0000000000000000100010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00004400000000000000000000000000) 
14'h05bc : LOC =         127'b0000000000000001000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00008400000000000000000000000000) 
14'h1561 : LOC =         127'b0000000000000010000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00010400000000000000000000000000) 
14'h34db : LOC =         127'b0000000000000100000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00020400000000000000000000000000) 
14'h34d8 : LOC =         127'b0000000000001000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00040400000000000000000000000000) 
14'h34de : LOC =         127'b0000000000010000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00080400000000000000000000000000) 
14'h34d2 : LOC =         127'b0000000000100000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00100400000000000000000000000000) 
14'h34ca : LOC =         127'b0000000001000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00200400000000000000000000000000) 
14'h34fa : LOC =         127'b0000000010000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00400400000000000000000000000000) 
14'h349a : LOC =         127'b0000000100000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00800400000000000000000000000000) 
14'h345a : LOC =         127'b0000001000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x01000400000000000000000000000000) 
14'h35da : LOC =         127'b0000010000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x02000400000000000000000000000000) 
14'h36da : LOC =         127'b0000100000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x04000400000000000000000000000000) 
14'h30da : LOC =         127'b0001000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x08000400000000000000000000000000) 
14'h3cda : LOC =         127'b0010000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x10000400000000000000000000000000) 
14'h24da : LOC =         127'b0100000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x20000400000000000000000000000000) 
14'h14da : LOC =         127'b1000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x40000400000000000000000000000000) 
14'h2ac3 : LOC =         127'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // S (0x00000800000000000000000000000000) 
14'h3c32 : LOC =         127'b0000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00001800000000000000000000000000) 
14'h0721 : LOC =         127'b0000000000000000010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00002800000000000000000000000000) 
14'h3270 : LOC =         127'b0000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00004800000000000000000000000000) 
14'h1ba5 : LOC =         127'b0000000000000001000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00008800000000000000000000000000) 
14'h0b78 : LOC =         127'b0000000000000010000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00010800000000000000000000000000) 
14'h2ac2 : LOC =         127'b0000000000000100000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00020800000000000000000000000000) 
14'h2ac1 : LOC =         127'b0000000000001000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00040800000000000000000000000000) 
14'h2ac7 : LOC =         127'b0000000000010000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00080800000000000000000000000000) 
14'h2acb : LOC =         127'b0000000000100000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00100800000000000000000000000000) 
14'h2ad3 : LOC =         127'b0000000001000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00200800000000000000000000000000) 
14'h2ae3 : LOC =         127'b0000000010000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00400800000000000000000000000000) 
14'h2a83 : LOC =         127'b0000000100000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00800800000000000000000000000000) 
14'h2a43 : LOC =         127'b0000001000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x01000800000000000000000000000000) 
14'h2bc3 : LOC =         127'b0000010000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x02000800000000000000000000000000) 
14'h28c3 : LOC =         127'b0000100000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x04000800000000000000000000000000) 
14'h2ec3 : LOC =         127'b0001000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x08000800000000000000000000000000) 
14'h22c3 : LOC =         127'b0010000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x10000800000000000000000000000000) 
14'h3ac3 : LOC =         127'b0100000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x20000800000000000000000000000000) 
14'h0ac3 : LOC =         127'b1000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x40000800000000000000000000000000) 
14'h16f1 : LOC =         127'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // S (0x00001000000000000000000000000000) 
14'h3b13 : LOC =         127'b0000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00003000000000000000000000000000) 
14'h0e42 : LOC =         127'b0000000000000000101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00005000000000000000000000000000) 
14'h2797 : LOC =         127'b0000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00009000000000000000000000000000) 
14'h374a : LOC =         127'b0000000000000010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00011000000000000000000000000000) 
14'h16f0 : LOC =         127'b0000000000000100001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00021000000000000000000000000000) 
14'h16f3 : LOC =         127'b0000000000001000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00041000000000000000000000000000) 
14'h16f5 : LOC =         127'b0000000000010000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00081000000000000000000000000000) 
14'h16f9 : LOC =         127'b0000000000100000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00101000000000000000000000000000) 
14'h16e1 : LOC =         127'b0000000001000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00201000000000000000000000000000) 
14'h16d1 : LOC =         127'b0000000010000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00401000000000000000000000000000) 
14'h16b1 : LOC =         127'b0000000100000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00801000000000000000000000000000) 
14'h1671 : LOC =         127'b0000001000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x01001000000000000000000000000000) 
14'h17f1 : LOC =         127'b0000010000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x02001000000000000000000000000000) 
14'h14f1 : LOC =         127'b0000100000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x04001000000000000000000000000000) 
14'h12f1 : LOC =         127'b0001000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x08001000000000000000000000000000) 
14'h1ef1 : LOC =         127'b0010000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x10001000000000000000000000000000) 
14'h06f1 : LOC =         127'b0100000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x20001000000000000000000000000000) 
14'h36f1 : LOC =         127'b1000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x40001000000000000000000000000000) 
14'h2de2 : LOC =         127'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // S (0x00002000000000000000000000000000) 
14'h3551 : LOC =         127'b0000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00006000000000000000000000000000) 
14'h1c84 : LOC =         127'b0000000000000001010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x0000a000000000000000000000000000) 
14'h0c59 : LOC =         127'b0000000000000010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00012000000000000000000000000000) 
14'h2de3 : LOC =         127'b0000000000000100010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00022000000000000000000000000000) 
14'h2de0 : LOC =         127'b0000000000001000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00042000000000000000000000000000) 
14'h2de6 : LOC =         127'b0000000000010000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00082000000000000000000000000000) 
14'h2dea : LOC =         127'b0000000000100000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00102000000000000000000000000000) 
14'h2df2 : LOC =         127'b0000000001000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00202000000000000000000000000000) 
14'h2dc2 : LOC =         127'b0000000010000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00402000000000000000000000000000) 
14'h2da2 : LOC =         127'b0000000100000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00802000000000000000000000000000) 
14'h2d62 : LOC =         127'b0000001000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x01002000000000000000000000000000) 
14'h2ce2 : LOC =         127'b0000010000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x02002000000000000000000000000000) 
14'h2fe2 : LOC =         127'b0000100000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x04002000000000000000000000000000) 
14'h29e2 : LOC =         127'b0001000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x08002000000000000000000000000000) 
14'h25e2 : LOC =         127'b0010000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x10002000000000000000000000000000) 
14'h3de2 : LOC =         127'b0100000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x20002000000000000000000000000000) 
14'h0de2 : LOC =         127'b1000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x40002000000000000000000000000000) 
14'h18b3 : LOC =         127'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // S (0x00004000000000000000000000000000) 
14'h29d5 : LOC =         127'b0000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x0000c000000000000000000000000000) 
14'h3908 : LOC =         127'b0000000000000010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00014000000000000000000000000000) 
14'h18b2 : LOC =         127'b0000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00024000000000000000000000000000) 
14'h18b1 : LOC =         127'b0000000000001000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00044000000000000000000000000000) 
14'h18b7 : LOC =         127'b0000000000010000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00084000000000000000000000000000) 
14'h18bb : LOC =         127'b0000000000100000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00104000000000000000000000000000) 
14'h18a3 : LOC =         127'b0000000001000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00204000000000000000000000000000) 
14'h1893 : LOC =         127'b0000000010000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00404000000000000000000000000000) 
14'h18f3 : LOC =         127'b0000000100000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00804000000000000000000000000000) 
14'h1833 : LOC =         127'b0000001000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x01004000000000000000000000000000) 
14'h19b3 : LOC =         127'b0000010000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x02004000000000000000000000000000) 
14'h1ab3 : LOC =         127'b0000100000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x04004000000000000000000000000000) 
14'h1cb3 : LOC =         127'b0001000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x08004000000000000000000000000000) 
14'h10b3 : LOC =         127'b0010000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x10004000000000000000000000000000) 
14'h08b3 : LOC =         127'b0100000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x20004000000000000000000000000000) 
14'h38b3 : LOC =         127'b1000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x40004000000000000000000000000000) 
14'h3166 : LOC =         127'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // S (0x00008000000000000000000000000000) 
14'h10dd : LOC =         127'b0000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00018000000000000000000000000000) 
14'h3167 : LOC =         127'b0000000000000101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00028000000000000000000000000000) 
14'h3164 : LOC =         127'b0000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00048000000000000000000000000000) 
14'h3162 : LOC =         127'b0000000000010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00088000000000000000000000000000) 
14'h316e : LOC =         127'b0000000000100001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00108000000000000000000000000000) 
14'h3176 : LOC =         127'b0000000001000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00208000000000000000000000000000) 
14'h3146 : LOC =         127'b0000000010000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00408000000000000000000000000000) 
14'h3126 : LOC =         127'b0000000100000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00808000000000000000000000000000) 
14'h31e6 : LOC =         127'b0000001000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x01008000000000000000000000000000) 
14'h3066 : LOC =         127'b0000010000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x02008000000000000000000000000000) 
14'h3366 : LOC =         127'b0000100000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x04008000000000000000000000000000) 
14'h3566 : LOC =         127'b0001000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x08008000000000000000000000000000) 
14'h3966 : LOC =         127'b0010000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x10008000000000000000000000000000) 
14'h2166 : LOC =         127'b0100000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x20008000000000000000000000000000) 
14'h1166 : LOC =         127'b1000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x40008000000000000000000000000000) 
14'h21bb : LOC =         127'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // S (0x00010000000000000000000000000000) 
14'h21ba : LOC =         127'b0000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00030000000000000000000000000000) 
14'h21b9 : LOC =         127'b0000000000001010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00050000000000000000000000000000) 
14'h21bf : LOC =         127'b0000000000010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00090000000000000000000000000000) 
14'h21b3 : LOC =         127'b0000000000100010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00110000000000000000000000000000) 
14'h21ab : LOC =         127'b0000000001000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00210000000000000000000000000000) 
14'h219b : LOC =         127'b0000000010000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00410000000000000000000000000000) 
14'h21fb : LOC =         127'b0000000100000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00810000000000000000000000000000) 
14'h213b : LOC =         127'b0000001000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x01010000000000000000000000000000) 
14'h20bb : LOC =         127'b0000010000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x02010000000000000000000000000000) 
14'h23bb : LOC =         127'b0000100000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x04010000000000000000000000000000) 
14'h25bb : LOC =         127'b0001000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x08010000000000000000000000000000) 
14'h29bb : LOC =         127'b0010000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x10010000000000000000000000000000) 
14'h31bb : LOC =         127'b0100000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x20010000000000000000000000000000) 
14'h01bb : LOC =         127'b1000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x40010000000000000000000000000000) 
14'h0001 : LOC =         127'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // S (0x00020000000000000000000000000000) 
14'h0003 : LOC =         127'b0000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00060000000000000000000000000000) 
14'h0005 : LOC =         127'b0000000000010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x000a0000000000000000000000000000) 
14'h0009 : LOC =         127'b0000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00120000000000000000000000000000) 
14'h0011 : LOC =         127'b0000000001000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00220000000000000000000000000000) 
14'h0021 : LOC =         127'b0000000010000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00420000000000000000000000000000) 
14'h0041 : LOC =         127'b0000000100000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00820000000000000000000000000000) 
14'h0081 : LOC =         127'b0000001000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x01020000000000000000000000000000) 
14'h0101 : LOC =         127'b0000010000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x02020000000000000000000000000000) 
14'h0201 : LOC =         127'b0000100000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x04020000000000000000000000000000) 
14'h0401 : LOC =         127'b0001000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x08020000000000000000000000000000) 
14'h0801 : LOC =         127'b0010000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x10020000000000000000000000000000) 
14'h1001 : LOC =         127'b0100000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x20020000000000000000000000000000) 
14'h2001 : LOC =         127'b1000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x40020000000000000000000000000000) 
14'h0002 : LOC =         127'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // S (0x00040000000000000000000000000000) 
14'h0006 : LOC =         127'b0000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x000c0000000000000000000000000000) 
14'h000a : LOC =         127'b0000000000101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00140000000000000000000000000000) 
14'h0012 : LOC =         127'b0000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00240000000000000000000000000000) 
14'h0022 : LOC =         127'b0000000010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00440000000000000000000000000000) 
14'h0042 : LOC =         127'b0000000100001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00840000000000000000000000000000) 
14'h0082 : LOC =         127'b0000001000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x01040000000000000000000000000000) 
14'h0102 : LOC =         127'b0000010000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x02040000000000000000000000000000) 
14'h0202 : LOC =         127'b0000100000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x04040000000000000000000000000000) 
14'h0402 : LOC =         127'b0001000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x08040000000000000000000000000000) 
14'h0802 : LOC =         127'b0010000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x10040000000000000000000000000000) 
14'h1002 : LOC =         127'b0100000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x20040000000000000000000000000000) 
14'h2002 : LOC =         127'b1000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x40040000000000000000000000000000) 
14'h0004 : LOC =         127'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // S (0x00080000000000000000000000000000) 
14'h000c : LOC =         127'b0000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00180000000000000000000000000000) 
14'h0014 : LOC =         127'b0000000001010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00280000000000000000000000000000) 
14'h0024 : LOC =         127'b0000000010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00480000000000000000000000000000) 
14'h0044 : LOC =         127'b0000000100010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00880000000000000000000000000000) 
14'h0084 : LOC =         127'b0000001000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x01080000000000000000000000000000) 
14'h0104 : LOC =         127'b0000010000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x02080000000000000000000000000000) 
14'h0204 : LOC =         127'b0000100000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x04080000000000000000000000000000) 
14'h0404 : LOC =         127'b0001000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x08080000000000000000000000000000) 
14'h0804 : LOC =         127'b0010000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x10080000000000000000000000000000) 
14'h1004 : LOC =         127'b0100000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x20080000000000000000000000000000) 
14'h2004 : LOC =         127'b1000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x40080000000000000000000000000000) 
14'h0008 : LOC =         127'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // S (0x00100000000000000000000000000000) 
14'h0018 : LOC =         127'b0000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00300000000000000000000000000000) 
14'h0028 : LOC =         127'b0000000010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00500000000000000000000000000000) 
14'h0048 : LOC =         127'b0000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00900000000000000000000000000000) 
14'h0088 : LOC =         127'b0000001000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x01100000000000000000000000000000) 
14'h0108 : LOC =         127'b0000010000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x02100000000000000000000000000000) 
14'h0208 : LOC =         127'b0000100000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x04100000000000000000000000000000) 
14'h0408 : LOC =         127'b0001000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x08100000000000000000000000000000) 
14'h0808 : LOC =         127'b0010000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x10100000000000000000000000000000) 
14'h1008 : LOC =         127'b0100000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x20100000000000000000000000000000) 
14'h2008 : LOC =         127'b1000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x40100000000000000000000000000000) 
14'h0010 : LOC =         127'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // S (0x00200000000000000000000000000000) 
14'h0030 : LOC =         127'b0000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00600000000000000000000000000000) 
14'h0050 : LOC =         127'b0000000101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00a00000000000000000000000000000) 
14'h0090 : LOC =         127'b0000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x01200000000000000000000000000000) 
14'h0110 : LOC =         127'b0000010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x02200000000000000000000000000000) 
14'h0210 : LOC =         127'b0000100001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x04200000000000000000000000000000) 
14'h0410 : LOC =         127'b0001000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x08200000000000000000000000000000) 
14'h0810 : LOC =         127'b0010000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x10200000000000000000000000000000) 
14'h1010 : LOC =         127'b0100000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x20200000000000000000000000000000) 
14'h2010 : LOC =         127'b1000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x40200000000000000000000000000000) 
14'h0020 : LOC =         127'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // S (0x00400000000000000000000000000000) 
14'h0060 : LOC =         127'b0000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x00c00000000000000000000000000000) 
14'h00a0 : LOC =         127'b0000001010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x01400000000000000000000000000000) 
14'h0120 : LOC =         127'b0000010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x02400000000000000000000000000000) 
14'h0220 : LOC =         127'b0000100010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x04400000000000000000000000000000) 
14'h0420 : LOC =         127'b0001000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x08400000000000000000000000000000) 
14'h0820 : LOC =         127'b0010000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x10400000000000000000000000000000) 
14'h1020 : LOC =         127'b0100000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x20400000000000000000000000000000) 
14'h2020 : LOC =         127'b1000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x40400000000000000000000000000000) 
14'h0040 : LOC =         127'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // S (0x00800000000000000000000000000000) 
14'h00c0 : LOC =         127'b0000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x01800000000000000000000000000000) 
14'h0140 : LOC =         127'b0000010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x02800000000000000000000000000000) 
14'h0240 : LOC =         127'b0000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x04800000000000000000000000000000) 
14'h0440 : LOC =         127'b0001000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x08800000000000000000000000000000) 
14'h0840 : LOC =         127'b0010000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x10800000000000000000000000000000) 
14'h1040 : LOC =         127'b0100000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x20800000000000000000000000000000) 
14'h2040 : LOC =         127'b1000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x40800000000000000000000000000000) 
14'h0080 : LOC =         127'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // S (0x01000000000000000000000000000000) 
14'h0180 : LOC =         127'b0000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x03000000000000000000000000000000) 
14'h0280 : LOC =         127'b0000101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x05000000000000000000000000000000) 
14'h0480 : LOC =         127'b0001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x09000000000000000000000000000000) 
14'h0880 : LOC =         127'b0010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x11000000000000000000000000000000) 
14'h1080 : LOC =         127'b0100001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x21000000000000000000000000000000) 
14'h2080 : LOC =         127'b1000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x41000000000000000000000000000000) 
14'h0100 : LOC =         127'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // S (0x02000000000000000000000000000000) 
14'h0300 : LOC =         127'b0000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x06000000000000000000000000000000) 
14'h0500 : LOC =         127'b0001010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x0a000000000000000000000000000000) 
14'h0900 : LOC =         127'b0010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x12000000000000000000000000000000) 
14'h1100 : LOC =         127'b0100010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x22000000000000000000000000000000) 
14'h2100 : LOC =         127'b1000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x42000000000000000000000000000000) 
14'h0200 : LOC =         127'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // S (0x04000000000000000000000000000000) 
14'h0600 : LOC =         127'b0001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x0c000000000000000000000000000000) 
14'h0a00 : LOC =         127'b0010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x14000000000000000000000000000000) 
14'h1200 : LOC =         127'b0100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x24000000000000000000000000000000) 
14'h2200 : LOC =         127'b1000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x44000000000000000000000000000000) 
14'h0400 : LOC =         127'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // S (0x08000000000000000000000000000000) 
14'h0c00 : LOC =         127'b0011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x18000000000000000000000000000000) 
14'h1400 : LOC =         127'b0101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x28000000000000000000000000000000) 
14'h2400 : LOC =         127'b1001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x48000000000000000000000000000000) 
14'h0800 : LOC =         127'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // S (0x10000000000000000000000000000000) 
14'h1800 : LOC =         127'b0110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x30000000000000000000000000000000) 
14'h2800 : LOC =         127'b1010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x50000000000000000000000000000000) 
14'h1000 : LOC =         127'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // S (0x20000000000000000000000000000000) 
14'h3000 : LOC =         127'b1100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // D (0x60000000000000000000000000000000) 
14'h2000 : LOC =         127'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // S (0x40000000000000000000000000000000) 
 
            default: LOC <= 0;
        endcase
        OUT <= LOC ^ IN;
    end
endmodule


module dec_top (input [140:0] IN, 
    output wire [126:0] OUT, 
    output reg [13:0] SYN, 
    output reg ERR, SGL, DBL,
    input clk 
);


    wire [13:0] CHK;
    assign CHK = IN[140:127];


    always @(*) begin
       SYN[0] <= CHK[0] ^ IN[0]^ IN[5]^ IN[6]^ IN[8]^ IN[9]^ IN[13]^ IN[14]^ IN[15]^ IN[17]^ IN[18]^ IN[19]^
              IN[22]^ IN[27]^ IN[28]^ IN[29]^ IN[30]^ IN[33]^ IN[34]^ IN[37]^ IN[39]^ IN[43]^
              IN[44]^ IN[45]^ IN[46]^ IN[48]^ IN[50]^ IN[51]^ IN[53]^ IN[57]^ IN[59]^ IN[61]^
              IN[64]^ IN[66]^ IN[68]^ IN[70]^ IN[72]^ IN[75]^ IN[77]^ IN[78]^ IN[80]^ IN[81]^
              IN[86]^ IN[88]^ IN[92]^ IN[93]^ IN[100]^ IN[101]^ IN[102]^ IN[103]^ IN[104]^ IN[105]^
              IN[107]^ IN[108]^ IN[110]^ IN[112]^ IN[113];

       SYN[1] <= CHK[1] ^ IN[0]^ IN[1]^ IN[5]^ IN[7]^ IN[8]^ IN[10]^ IN[13]^ IN[16]^ IN[17]^ IN[20]^ IN[22]^
              IN[23]^ IN[27]^ IN[31]^ IN[33]^ IN[35]^ IN[37]^ IN[38]^ IN[39]^ IN[40]^ IN[43]^
              IN[47]^ IN[48]^ IN[49]^ IN[50]^ IN[52]^ IN[53]^ IN[54]^ IN[57]^ IN[58]^ IN[59]^
              IN[60]^ IN[61]^ IN[62]^ IN[64]^ IN[65]^ IN[66]^ IN[67]^ IN[68]^ IN[69]^ IN[70]^
              IN[71]^ IN[72]^ IN[73]^ IN[75]^ IN[76]^ IN[77]^ IN[79]^ IN[80]^ IN[82]^ IN[86]^
              IN[87]^ IN[88]^ IN[89]^ IN[92]^ IN[94]^ IN[100]^ IN[106]^ IN[107]^ IN[109]^ IN[110]^
              IN[111]^ IN[112]^ IN[114];

       SYN[2] <= CHK[2] ^  IN[0]^ IN[1]^ IN[2]^ IN[5]^ IN[11]^ IN[13]^ IN[15]^ IN[19]^ IN[21]^ IN[22]^ IN[23]^
               IN[24]^ IN[27]^ IN[29]^ IN[30]^ IN[32]^ IN[33]^ IN[36]^ IN[37]^ IN[38]^ IN[40]^
               IN[41]^ IN[43]^ IN[45]^ IN[46]^ IN[49]^ IN[54]^ IN[55]^ IN[57]^ IN[58]^ IN[60]^
               IN[62]^ IN[63]^ IN[64]^ IN[65]^ IN[67]^ IN[69]^ IN[71]^ IN[73]^ IN[74]^ IN[75]^
               IN[76]^ IN[83]^ IN[86]^ IN[87]^ IN[89]^ IN[90]^ IN[92]^ IN[95]^ IN[100]^ IN[102]^
               IN[103]^ IN[104]^ IN[105]^ IN[111]^ IN[115];

       SYN[3] <= CHK[3] ^  IN[1]^ IN[2]^ IN[3]^ IN[6]^ IN[12]^ IN[14]^ IN[16]^ IN[20]^ IN[22]^ IN[23]^ IN[24]^
               IN[25]^ IN[28]^ IN[30]^ IN[31]^ IN[33]^ IN[34]^ IN[37]^ IN[38]^ IN[39]^ IN[41]^ IN[42]^
               IN[44]^ IN[46]^ IN[47]^ IN[50]^ IN[55]^ IN[56]^ IN[58]^ IN[59]^ IN[61]^ IN[63]^ IN[64]^
               IN[65]^ IN[66]^ IN[68]^ IN[70]^ IN[72]^ IN[74]^ IN[75]^ IN[76]^ IN[77]^ IN[84]^ IN[87]^
               IN[88]^ IN[90]^ IN[91]^ IN[93]^ IN[96]^ IN[101]^ IN[103]^ IN[104]^ IN[105]^ IN[106]^
               IN[112]^ IN[116];

       SYN[4] <= CHK[4] ^  IN[0]^ IN[2]^ IN[3]^ IN[4]^ IN[5]^ IN[6]^ IN[7]^ IN[8]^ IN[9]^ IN[14]^ IN[18]^ IN[19]^
               IN[21]^ IN[22]^ IN[23]^ IN[24]^ IN[25]^ IN[26]^ IN[27]^ IN[28]^ IN[30]^ IN[31]^ IN[32]^
               IN[33]^ IN[35]^ IN[37]^ IN[38]^ IN[40]^ IN[42]^ IN[44]^ IN[46]^ IN[47]^ IN[50]^ IN[53]^
               IN[56]^ IN[60]^ IN[61]^ IN[62]^ IN[65]^ IN[67]^ IN[68]^ IN[69]^ IN[70]^ IN[71]^ IN[72]^
               IN[73]^ IN[76]^ IN[80]^ IN[81]^ IN[85]^ IN[86]^ IN[89]^ IN[91]^ IN[93]^ IN[94]^ IN[97]^
               IN[100]^ IN[101]^ IN[103]^ IN[106]^ IN[108]^ IN[110]^ IN[112]^ IN[117];

       SYN[5] <= CHK[5] ^  IN[0]^ IN[1]^ IN[3]^ IN[4]^ IN[7]^ IN[10]^ IN[13]^ IN[14]^ IN[17]^ IN[18]^ IN[20]^ IN[23]^
               IN[24]^ IN[25]^ IN[26]^ IN[30]^ IN[31]^ IN[32]^ IN[36]^ IN[37]^ IN[38]^ IN[41]^ IN[44]^																		   
               IN[46]^ IN[47]^ IN[50]^ IN[53]^ IN[54]^ IN[59]^ IN[62]^ IN[63]^ IN[64]^ IN[69]^ IN[71]^
               IN[73]^ IN[74]^ IN[75]^ IN[78]^ IN[80]^ IN[82]^ IN[87]^ IN[88]^ IN[90]^ IN[93]^ IN[94]^
               IN[95]^ IN[98]^ IN[100]^ IN[103]^ IN[105]^ IN[108]^ IN[109]^ IN[110]^ IN[111]^ IN[112]^
               IN[118];

       SYN[6] <= CHK[6] ^  IN[0]^ IN[1]^ IN[2]^ IN[4]^ IN[6]^ IN[9]^ IN[11]^ IN[13]^ IN[17]^ IN[21]^ IN[22]^ IN[24]^
               IN[25]^ IN[26]^ IN[28]^ IN[29]^ IN[30]^ IN[31]^ IN[32]^ IN[34]^ IN[38]^ IN[42]^ IN[43]^
               IN[44]^ IN[46]^ IN[47]^ IN[50]^ IN[53]^ IN[54]^ IN[55]^ IN[57]^ IN[59]^ IN[60]^ IN[61]^
               IN[63]^ IN[65]^ IN[66]^ IN[68]^ IN[74]^ IN[76]^ IN[77]^ IN[78]^ IN[79]^ IN[80]^ IN[83]^
               IN[86]^ IN[89]^ IN[91]^ IN[92]^ IN[93]^ IN[94]^ IN[95]^ IN[96]^ IN[99]^ IN[100]^ IN[102]^
               IN[103]^ IN[105]^ IN[106]^ IN[107]^ IN[108]^ IN[109]^ IN[111]^ IN[119];

       SYN[7] <= CHK[7] ^  IN[1]^ IN[2]^ IN[3]^ IN[5]^ IN[7]^ IN[10]^ IN[12]^ IN[14]^ IN[18]^ IN[22]^ IN[23]^ IN[25]^
               IN[26]^ IN[27]^ IN[29]^ IN[30]^ IN[31]^ IN[32]^ IN[33]^ IN[35]^ IN[39]^ IN[43]^ IN[44]^
               IN[45]^ IN[47]^ IN[48]^ IN[51]^ IN[54]^ IN[55]^ IN[56]^ IN[58]^ IN[60]^ IN[61]^ IN[62]^
               IN[64]^ IN[66]^ IN[67]^ IN[69]^ IN[75]^ IN[77]^ IN[78]^ IN[79]^ IN[80]^ IN[81]^ IN[84]^ 
               IN[87]^ IN[90]^ IN[92]^ IN[93]^ IN[94]^ IN[95]^ IN[96]^ IN[97]^ IN[100]^ IN[101]^ IN[103]^
               IN[104]^ IN[106]^ IN[107]^ IN[108]^ IN[109]^ IN[110]^ IN[112]^ IN[120];

       SYN[8] <= CHK[8] ^  IN[0]^ IN[2]^ IN[3]^ IN[4]^ IN[5]^ IN[9]^ IN[11]^ IN[14]^ IN[17]^ IN[18]^ IN[22]^ IN[23]^
               IN[24]^ IN[26]^ IN[29]^ IN[31]^ IN[32]^ IN[36]^ IN[37]^ IN[39]^ IN[40]^ IN[43]^ IN[49]^
               IN[50]^ IN[51]^ IN[52]^ IN[53]^ IN[55]^ IN[56]^ IN[62]^ IN[63]^ IN[64]^ IN[65]^ IN[66]^
               IN[67]^ IN[72]^ IN[75]^ IN[76]^ IN[77]^ IN[79]^ IN[82]^ IN[85]^ IN[86]^ IN[91]^ IN[92]^
               IN[94]^ IN[95]^ IN[96]^ IN[97]^ IN[98]^ IN[100]^ IN[103]^ IN[109]^ IN[111]^ IN[112]^ IN[121];

       SYN[9] <= CHK[9] ^  IN[0]^ IN[1]^ IN[3]^ IN[4]^ IN[8]^ IN[9]^ IN[10]^ IN[12]^ IN[13]^ IN[14]^ IN[17]^ IN[22]^ IN[23]^
               IN[24]^ IN[25]^ IN[28]^ IN[29]^ IN[32]^ IN[34]^ IN[38]^ IN[39]^ IN[40]^ IN[41]^ IN[43]^ IN[45]^
               IN[46]^ IN[48]^ IN[52]^ IN[54]^ IN[56]^ IN[59]^ IN[61]^ IN[63]^ IN[65]^ IN[67]^ IN[70]^ IN[72]^
               IN[73]^ IN[75]^ IN[76]^ IN[81]^ IN[83]^ IN[87]^ IN[88]^ IN[95]^ IN[96]^ IN[97]^ IN[98]^ IN[99]^
               IN[100]^ IN[102]^ IN[103]^ IN[105]^ IN[107]^ IN[108]^ IN[122];

       SYN[10] <= CHK[10] ^ IN[1]^ IN[2]^ IN[4]^ IN[5]^ IN[9]^ IN[10]^ IN[11]^ IN[13]^ IN[14]^ IN[15]^ IN[18]^ IN[23]^ IN[24]^
               IN[25]^ IN[26]^ IN[29]^ IN[30]^ IN[33]^ IN[35]^ IN[39]^ IN[40]^ IN[41]^ IN[42]^ IN[44]^ IN[46]^
               IN[47]^ IN[49]^ IN[53]^ IN[55]^ IN[57]^ IN[60]^ IN[62]^ IN[64]^ IN[66]^ IN[68]^ IN[71]^ IN[73]^
               IN[74]^ IN[76]^ IN[77]^ IN[82]^ IN[84]^ IN[88]^ IN[89]^ IN[96]^ IN[97]^ IN[98]^ IN[99]^ IN[100]^ 
               IN[101]^ IN[103]^ IN[104]^ IN[106]^ IN[108]^ IN[109]^ IN[123];

       SYN[11] <= CHK[11] ^ IN[2]^ IN[3]^ IN[5]^ IN[6]^ IN[10]^ IN[11]^ IN[12]^ IN[14]^ IN[15]^ IN[16]^ IN[19]^ IN[24]^ IN[25]^
               IN[26]^ IN[27]^ IN[30]^ IN[31]^ IN[34]^ IN[36]^ IN[40]^ IN[41]^ IN[42]^ IN[43]^ IN[45]^ IN[47]^ IN[48]^
               IN[50]^ IN[54]^ IN[56]^ IN[58]^ IN[61]^ IN[63]^ IN[65]^ IN[67]^ IN[69]^ IN[72]^ IN[74]^ IN[75]^ IN[77]^
               IN[78]^ IN[83]^ IN[85]^ IN[89]^ IN[90]^ IN[97]^ IN[98]^ IN[99]^ IN[100]^ IN[101]^ IN[102]^ IN[104]^
               IN[105]^ IN[107]^ IN[109]^ IN[110]^ IN[124];

       SYN[12] <= CHK[12] ^ IN[3]^ IN[4]^ IN[6]^ IN[7]^ IN[11]^ IN[12]^IN[13]^ IN[15]^ IN[16]^ IN[17]^ IN[20]^ IN[25]^ IN[26]^
               IN[27]^ IN[28]^ IN[31]^ IN[32]^ IN[35]^ IN[37]^ IN[41]^ IN[42]^ IN[43]^ IN[44]^ IN[46]^ IN[48]^
               IN[49]^ IN[51]^ IN[55]^ IN[57]^ IN[59]^ IN[62]^ IN[64]^ IN[66]^ IN[68]^ IN[70]^ IN[73]^ IN[75]^
               IN[76]^ IN[78]^ IN[79]^ IN[84]^ IN[86]^ IN[90]^ IN[91]^ IN[98]^ IN[99]^ IN[100]^ IN[101]^ IN[102]^
               IN[103]^ IN[105]^ IN[106]^ IN[108]^ IN[110]^ IN[111]^ IN[125];

       SYN[13] <= CHK[13] ^  IN[4]^ IN[5]^ IN[7]^ IN[8]^ IN[12]^ IN[13]^ IN[14]^ IN[16]^ IN[17]^ IN[18]^ IN[21]^ IN[26]^ IN[27]^
                IN[28]^ IN[29]^ IN[32]^ IN[33]^ IN[36]^ IN[38]^ IN[42]^ IN[43]^ IN[44]^ IN[45]^ IN[47]^ IN[49]^
                IN[50]^ IN[52]^ IN[56]^ IN[58]^ IN[60]^ IN[63]^ IN[65]^ IN[67]^ IN[69]^ IN[71]^ IN[74]^ IN[76]^
                IN[77]^ IN[79]^ IN[80]^ IN[85]^ IN[87]^ IN[91]^ IN[92]^ IN[99]^ IN[100]^ IN[101]^ IN[102]^
                IN[103]^ IN[104]^ IN[106]^ IN[107]^ IN[109]^ IN[111]^ IN[112]^ IN[126];


      
        ERR <= |SYN;
        SGL <= ^SYN & ERR;
        DBL <= ~^SYN & ERR;
    end

corrector corr_mod (.IN(IN[126:0]), .SYN(SYN), .OUT(OUT));
    
endmodule



