//
// decoder for Hsiaod 64 bit DEC
//
// Authors: Joseph Crowe and Matt Markwell
//


module corrector (input [62:0] IN, 
    input [11:0] SYN,
    output reg [62:0] OUT
);

reg [62:0] LOC;

    always @(*) begin
        case(SYN)

    12'h539 : LOC <=          63'b000000000000000000000000000000000000000000000000000000000000001; // S (0x0000000000000001) 
//    12'hf4b : LOC <=          63'b000000000000000000000000000000000000000000000000000000000000011; // D (0x0000000000000003) 
//    12'h4e4 : LOC <=          63'b000000000000000000000000000000000000000000000000000000000000101; // D (0x0000000000000005) 
//    12'h683 : LOC <=          63'b000000000000000000000000000000000000000000000000000000000001001; // D (0x0000000000000009) 
//    12'h24d : LOC <=          63'b000000000000000000000000000000000000000000000000000000000010001; // D (0x0000000000000011) 
//    12'hbd1 : LOC <=          63'b000000000000000000000000000000000000000000000000000000000100001; // D (0x0000000000000021) 
//    12'hdd0 : LOC <=          63'b000000000000000000000000000000000000000000000000000000001000001; // D (0x0000000000000041) 
//    12'h1d2 : LOC <=          63'b000000000000000000000000000000000000000000000000000000010000001; // D (0x0000000000000081) 
//    12'hcef : LOC <=          63'b000000000000000000000000000000000000000000000000000000100000001; // D (0x0000000000000101) 
//    12'h3ac : LOC <=          63'b000000000000000000000000000000000000000000000000000001000000001; // D (0x0000000000000201) 
//    12'h813 : LOC <=          63'b000000000000000000000000000000000000000000000000000010000000001; // D (0x0000000000000401) 
//    12'ha54 : LOC <=          63'b000000000000000000000000000000000000000000000000000100000000001; // D (0x0000000000000801) 
//    12'heda : LOC <=          63'b000000000000000000000000000000000000000000000000001000000000001; // D (0x0000000000001001) 
//    12'h7c6 : LOC <=          63'b000000000000000000000000000000000000000000000000010000000000001; // D (0x0000000000002001) 
//    12'h0c7 : LOC <=          63'b000000000000000000000000000000000000000000000000100000000000001; // D (0x0000000000004001) 
//    12'hec5 : LOC <=          63'b000000000000000000000000000000000000000000000001000000000000001; // D (0x0000000000008001) 
//    12'h7f8 : LOC <=          63'b000000000000000000000000000000000000000000000010000000000000001; // D (0x0000000000010001) 
//    12'h0bb : LOC <=          63'b000000000000000000000000000000000000000000000100000000000000001; // D (0x0000000000020001) 
//    12'he3d : LOC <=          63'b000000000000000000000000000000000000000000001000000000000000001; // D (0x0000000000040001) 
//    12'h608 : LOC <=          63'b000000000000000000000000000000000000000000010000000000000000001; // D (0x0000000000080001) 
//    12'h35b : LOC <=          63'b000000000000000000000000000000000000000000100000000000000000001; // D (0x0000000000100001) 
//    12'h9fd : LOC <=          63'b000000000000000000000000000000000000000001000000000000000000001; // D (0x0000000000200001) 
//    12'h988 : LOC <=          63'b000000000000000000000000000000000000000010000000000000000000001; // D (0x0000000000400001) 
//    12'h962 : LOC <=          63'b000000000000000000000000000000000000000100000000000000000000001; // D (0x0000000000800001) 
//    12'h8b6 : LOC <=          63'b000000000000000000000000000000000000001000000000000000000000001; // D (0x0000000001000001) 
//    12'hb1e : LOC <=          63'b000000000000000000000000000000000000010000000000000000000000001; // D (0x0000000002000001) 
//    12'hc4e : LOC <=          63'b000000000000000000000000000000000000100000000000000000000000001; // D (0x0000000004000001) 
//    12'h2ee : LOC <=          63'b000000000000000000000000000000000001000000000000000000000000001; // D (0x0000000008000001) 
//    12'ha97 : LOC <=          63'b000000000000000000000000000000000010000000000000000000000000001; // D (0x0000000010000001) 
//    12'hf5c : LOC <=          63'b000000000000000000000000000000000100000000000000000000000000001; // D (0x0000000020000001) 
//    12'h4ca : LOC <=          63'b000000000000000000000000000000001000000000000000000000000000001; // D (0x0000000040000001) 
//    12'h6df : LOC <=          63'b000000000000000000000000000000010000000000000000000000000000001; // D (0x0000000080000001) 
//    12'h2f5 : LOC <=          63'b000000000000000000000000000000100000000000000000000000000000001; // D (0x0000000100000001) 
//    12'haa1 : LOC <=          63'b000000000000000000000000000001000000000000000000000000000000001; // D (0x0000000200000001) 
//    12'hf30 : LOC <=          63'b000000000000000000000000000010000000000000000000000000000000001; // D (0x0000000400000001) 
//    12'h412 : LOC <=          63'b000000000000000000000000000100000000000000000000000000000000001; // D (0x0000000800000001) 
//    12'h76f : LOC <=          63'b000000000000000000000000001000000000000000000000000000000000001; // D (0x0000001000000001) 
//    12'h195 : LOC <=          63'b000000000000000000000000010000000000000000000000000000000000001; // D (0x0000002000000001) 
//    12'hc61 : LOC <=          63'b000000000000000000000000100000000000000000000000000000000000001; // D (0x0000004000000001) 
//    12'h2b0 : LOC <=          63'b000000000000000000000001000000000000000000000000000000000000001; // D (0x0000008000000001) 
//    12'ha2b : LOC <=          63'b000000000000000000000010000000000000000000000000000000000000001; // D (0x0000010000000001) 
//    12'he24 : LOC <=          63'b000000000000000000000100000000000000000000000000000000000000001; // D (0x0000020000000001) 
//    12'h63a : LOC <=          63'b000000000000000000001000000000000000000000000000000000000000001; // D (0x0000040000000001) 
//    12'h33f : LOC <=          63'b000000000000000000010000000000000000000000000000000000000000001; // D (0x0000080000000001) 
//    12'h935 : LOC <=          63'b000000000000000000100000000000000000000000000000000000000000001; // D (0x0000100000000001) 
//    12'h818 : LOC <=          63'b000000000000000001000000000000000000000000000000000000000000001; // D (0x0000200000000001) 
//    12'ha42 : LOC <=          63'b000000000000000010000000000000000000000000000000000000000000001; // D (0x0000400000000001) 
//    12'hef6 : LOC <=          63'b000000000000000100000000000000000000000000000000000000000000001; // D (0x0000800000000001) 
//    12'h79e : LOC <=          63'b000000000000001000000000000000000000000000000000000000000000001; // D (0x0001000000000001) 
//    12'h077 : LOC <=          63'b000000000000010000000000000000000000000000000000000000000000001; // D (0x0002000000000001) 
//    12'hfa5 : LOC <=          63'b000000000000100000000000000000000000000000000000000000000000001; // D (0x0004000000000001) 
//    12'h538 : LOC <=          63'b000000000001000000000000000000000000000000000000000000000000001; // D (0x0008000000000001) 
//    12'h53b : LOC <=          63'b000000000010000000000000000000000000000000000000000000000000001; // D (0x0010000000000001) 
//    12'h53d : LOC <=          63'b000000000100000000000000000000000000000000000000000000000000001; // D (0x0020000000000001) 
//    12'h531 : LOC <=          63'b000000001000000000000000000000000000000000000000000000000000001; // D (0x0040000000000001) 
//    12'h529 : LOC <=          63'b000000010000000000000000000000000000000000000000000000000000001; // D (0x0080000000000001) 
//    12'h519 : LOC <=          63'b000000100000000000000000000000000000000000000000000000000000001; // D (0x0100000000000001) 
//    12'h579 : LOC <=          63'b000001000000000000000000000000000000000000000000000000000000001; // D (0x0200000000000001) 
//    12'h5b9 : LOC <=          63'b000010000000000000000000000000000000000000000000000000000000001; // D (0x0400000000000001) 
//    12'h439 : LOC <=          63'b000100000000000000000000000000000000000000000000000000000000001; // D (0x0800000000000001) 
//    12'h739 : LOC <=          63'b001000000000000000000000000000000000000000000000000000000000001; // D (0x1000000000000001) 
//    12'h139 : LOC <=          63'b010000000000000000000000000000000000000000000000000000000000001; // D (0x2000000000000001) 
//    12'hd39 : LOC <=          63'b100000000000000000000000000000000000000000000000000000000000001; // D (0x4000000000000001) 
    12'hf4b : LOC <=          63'b000000000000000000000000000000000000000000000000000000000000011; // D (0x0000000000000003) 
    12'ha72 : LOC <=          63'b000000000000000000000000000000000000000000000000000000000000010; // S (0x0000000000000002) 
//    12'hbaf : LOC <=          63'b000000000000000000000000000000000000000000000000000000000000110; // D (0x0000000000000006) 
//    12'h9c8 : LOC <=          63'b000000000000000000000000000000000000000000000000000000000001010; // D (0x000000000000000a) 
//    12'hd06 : LOC <=          63'b000000000000000000000000000000000000000000000000000000000010010; // D (0x0000000000000012) 
//    12'h49a : LOC <=          63'b000000000000000000000000000000000000000000000000000000000100010; // D (0x0000000000000022) 
//    12'h29b : LOC <=          63'b000000000000000000000000000000000000000000000000000000001000010; // D (0x0000000000000042) 
//    12'he99 : LOC <=          63'b000000000000000000000000000000000000000000000000000000010000010; // D (0x0000000000000082) 
//    12'h3a4 : LOC <=          63'b000000000000000000000000000000000000000000000000000000100000010; // D (0x0000000000000102) 
//    12'hce7 : LOC <=          63'b000000000000000000000000000000000000000000000000000001000000010; // D (0x0000000000000202) 
//    12'h758 : LOC <=          63'b000000000000000000000000000000000000000000000000000010000000010; // D (0x0000000000000402) 
//    12'h51f : LOC <=          63'b000000000000000000000000000000000000000000000000000100000000010; // D (0x0000000000000802) 
//    12'h191 : LOC <=          63'b000000000000000000000000000000000000000000000000001000000000010; // D (0x0000000000001002) 
//    12'h88d : LOC <=          63'b000000000000000000000000000000000000000000000000010000000000010; // D (0x0000000000002002) 
//    12'hf8c : LOC <=          63'b000000000000000000000000000000000000000000000000100000000000010; // D (0x0000000000004002) 
//    12'h18e : LOC <=          63'b000000000000000000000000000000000000000000000001000000000000010; // D (0x0000000000008002) 
//    12'h8b3 : LOC <=          63'b000000000000000000000000000000000000000000000010000000000000010; // D (0x0000000000010002) 
//    12'hff0 : LOC <=          63'b000000000000000000000000000000000000000000000100000000000000010; // D (0x0000000000020002) 
//    12'h176 : LOC <=          63'b000000000000000000000000000000000000000000001000000000000000010; // D (0x0000000000040002) 
//    12'h943 : LOC <=          63'b000000000000000000000000000000000000000000010000000000000000010; // D (0x0000000000080002) 
//    12'hc10 : LOC <=          63'b000000000000000000000000000000000000000000100000000000000000010; // D (0x0000000000100002) 
//    12'h6b6 : LOC <=          63'b000000000000000000000000000000000000000001000000000000000000010; // D (0x0000000000200002) 
//    12'h6c3 : LOC <=          63'b000000000000000000000000000000000000000010000000000000000000010; // D (0x0000000000400002) 
//    12'h629 : LOC <=          63'b000000000000000000000000000000000000000100000000000000000000010; // D (0x0000000000800002) 
//    12'h7fd : LOC <=          63'b000000000000000000000000000000000000001000000000000000000000010; // D (0x0000000001000002) 
//    12'h455 : LOC <=          63'b000000000000000000000000000000000000010000000000000000000000010; // D (0x0000000002000002) 
//    12'h305 : LOC <=          63'b000000000000000000000000000000000000100000000000000000000000010; // D (0x0000000004000002) 
//    12'hda5 : LOC <=          63'b000000000000000000000000000000000001000000000000000000000000010; // D (0x0000000008000002) 
//    12'h5dc : LOC <=          63'b000000000000000000000000000000000010000000000000000000000000010; // D (0x0000000010000002) 
//    12'h017 : LOC <=          63'b000000000000000000000000000000000100000000000000000000000000010; // D (0x0000000020000002) 
//    12'hb81 : LOC <=          63'b000000000000000000000000000000001000000000000000000000000000010; // D (0x0000000040000002) 
//    12'h994 : LOC <=          63'b000000000000000000000000000000010000000000000000000000000000010; // D (0x0000000080000002) 
//    12'hdbe : LOC <=          63'b000000000000000000000000000000100000000000000000000000000000010; // D (0x0000000100000002) 
//    12'h5ea : LOC <=          63'b000000000000000000000000000001000000000000000000000000000000010; // D (0x0000000200000002) 
//    12'h07b : LOC <=          63'b000000000000000000000000000010000000000000000000000000000000010; // D (0x0000000400000002) 
//    12'hb59 : LOC <=          63'b000000000000000000000000000100000000000000000000000000000000010; // D (0x0000000800000002) 
//    12'h824 : LOC <=          63'b000000000000000000000000001000000000000000000000000000000000010; // D (0x0000001000000002) 
//    12'hede : LOC <=          63'b000000000000000000000000010000000000000000000000000000000000010; // D (0x0000002000000002) 
//    12'h32a : LOC <=          63'b000000000000000000000000100000000000000000000000000000000000010; // D (0x0000004000000002) 
//    12'hdfb : LOC <=          63'b000000000000000000000001000000000000000000000000000000000000010; // D (0x0000008000000002) 
//    12'h560 : LOC <=          63'b000000000000000000000010000000000000000000000000000000000000010; // D (0x0000010000000002) 
//    12'h16f : LOC <=          63'b000000000000000000000100000000000000000000000000000000000000010; // D (0x0000020000000002) 
//    12'h971 : LOC <=          63'b000000000000000000001000000000000000000000000000000000000000010; // D (0x0000040000000002) 
//    12'hc74 : LOC <=          63'b000000000000000000010000000000000000000000000000000000000000010; // D (0x0000080000000002) 
//    12'h67e : LOC <=          63'b000000000000000000100000000000000000000000000000000000000000010; // D (0x0000100000000002) 
//    12'h753 : LOC <=          63'b000000000000000001000000000000000000000000000000000000000000010; // D (0x0000200000000002) 
//    12'h509 : LOC <=          63'b000000000000000010000000000000000000000000000000000000000000010; // D (0x0000400000000002) 
//    12'h1bd : LOC <=          63'b000000000000000100000000000000000000000000000000000000000000010; // D (0x0000800000000002) 
//    12'h8d5 : LOC <=          63'b000000000000001000000000000000000000000000000000000000000000010; // D (0x0001000000000002) 
//    12'hf3c : LOC <=          63'b000000000000010000000000000000000000000000000000000000000000010; // D (0x0002000000000002) 
//    12'h0ee : LOC <=          63'b000000000000100000000000000000000000000000000000000000000000010; // D (0x0004000000000002) 
//    12'ha73 : LOC <=          63'b000000000001000000000000000000000000000000000000000000000000010; // D (0x0008000000000002) 
//    12'ha70 : LOC <=          63'b000000000010000000000000000000000000000000000000000000000000010; // D (0x0010000000000002) 
//    12'ha76 : LOC <=          63'b000000000100000000000000000000000000000000000000000000000000010; // D (0x0020000000000002) 
//    12'ha7a : LOC <=          63'b000000001000000000000000000000000000000000000000000000000000010; // D (0x0040000000000002) 
//    12'ha62 : LOC <=          63'b000000010000000000000000000000000000000000000000000000000000010; // D (0x0080000000000002) 
//    12'ha52 : LOC <=          63'b000000100000000000000000000000000000000000000000000000000000010; // D (0x0100000000000002) 
//    12'ha32 : LOC <=          63'b000001000000000000000000000000000000000000000000000000000000010; // D (0x0200000000000002) 
//    12'haf2 : LOC <=          63'b000010000000000000000000000000000000000000000000000000000000010; // D (0x0400000000000002) 
//    12'hb72 : LOC <=          63'b000100000000000000000000000000000000000000000000000000000000010; // D (0x0800000000000002) 
//    12'h872 : LOC <=          63'b001000000000000000000000000000000000000000000000000000000000010; // D (0x1000000000000002) 
//    12'he72 : LOC <=          63'b010000000000000000000000000000000000000000000000000000000000010; // D (0x2000000000000002) 
//    12'h272 : LOC <=          63'b100000000000000000000000000000000000000000000000000000000000010; // D (0x4000000000000002) 
    12'h4e4 : LOC <=          63'b000000000000000000000000000000000000000000000000000000000000101; // D (0x0000000000000005) 
    12'hbaf : LOC <=          63'b000000000000000000000000000000000000000000000000000000000000110; // D (0x0000000000000006) 
    12'h1dd : LOC <=          63'b000000000000000000000000000000000000000000000000000000000000100; // S (0x0000000000000004) 
//    12'h267 : LOC <=          63'b000000000000000000000000000000000000000000000000000000000001100; // D (0x000000000000000c) 
//    12'h6a9 : LOC <=          63'b000000000000000000000000000000000000000000000000000000000010100; // D (0x0000000000000014) 
//    12'hf35 : LOC <=          63'b000000000000000000000000000000000000000000000000000000000100100; // D (0x0000000000000024) 
//    12'h934 : LOC <=          63'b000000000000000000000000000000000000000000000000000000001000100; // D (0x0000000000000044) 
//    12'h536 : LOC <=          63'b000000000000000000000000000000000000000000000000000000010000100; // D (0x0000000000000084) 
//    12'h80b : LOC <=          63'b000000000000000000000000000000000000000000000000000000100000100; // D (0x0000000000000104) 
//    12'h748 : LOC <=          63'b000000000000000000000000000000000000000000000000000001000000100; // D (0x0000000000000204) 
//    12'hcf7 : LOC <=          63'b000000000000000000000000000000000000000000000000000010000000100; // D (0x0000000000000404) 
//    12'heb0 : LOC <=          63'b000000000000000000000000000000000000000000000000000100000000100; // D (0x0000000000000804) 
//    12'ha3e : LOC <=          63'b000000000000000000000000000000000000000000000000001000000000100; // D (0x0000000000001004) 
//    12'h322 : LOC <=          63'b000000000000000000000000000000000000000000000000010000000000100; // D (0x0000000000002004) 
//    12'h423 : LOC <=          63'b000000000000000000000000000000000000000000000000100000000000100; // D (0x0000000000004004) 
//    12'ha21 : LOC <=          63'b000000000000000000000000000000000000000000000001000000000000100; // D (0x0000000000008004) 
//    12'h31c : LOC <=          63'b000000000000000000000000000000000000000000000010000000000000100; // D (0x0000000000010004) 
//    12'h45f : LOC <=          63'b000000000000000000000000000000000000000000000100000000000000100; // D (0x0000000000020004) 
//    12'had9 : LOC <=          63'b000000000000000000000000000000000000000000001000000000000000100; // D (0x0000000000040004) 
//    12'h2ec : LOC <=          63'b000000000000000000000000000000000000000000010000000000000000100; // D (0x0000000000080004) 
//    12'h7bf : LOC <=          63'b000000000000000000000000000000000000000000100000000000000000100; // D (0x0000000000100004) 
//    12'hd19 : LOC <=          63'b000000000000000000000000000000000000000001000000000000000000100; // D (0x0000000000200004) 
//    12'hd6c : LOC <=          63'b000000000000000000000000000000000000000010000000000000000000100; // D (0x0000000000400004) 
//    12'hd86 : LOC <=          63'b000000000000000000000000000000000000000100000000000000000000100; // D (0x0000000000800004) 
//    12'hc52 : LOC <=          63'b000000000000000000000000000000000000001000000000000000000000100; // D (0x0000000001000004) 
//    12'hffa : LOC <=          63'b000000000000000000000000000000000000010000000000000000000000100; // D (0x0000000002000004) 
//    12'h8aa : LOC <=          63'b000000000000000000000000000000000000100000000000000000000000100; // D (0x0000000004000004) 
//    12'h60a : LOC <=          63'b000000000000000000000000000000000001000000000000000000000000100; // D (0x0000000008000004) 
//    12'he73 : LOC <=          63'b000000000000000000000000000000000010000000000000000000000000100; // D (0x0000000010000004) 
//    12'hbb8 : LOC <=          63'b000000000000000000000000000000000100000000000000000000000000100; // D (0x0000000020000004) 
//    12'h02e : LOC <=          63'b000000000000000000000000000000001000000000000000000000000000100; // D (0x0000000040000004) 
//    12'h23b : LOC <=          63'b000000000000000000000000000000010000000000000000000000000000100; // D (0x0000000080000004) 
//    12'h611 : LOC <=          63'b000000000000000000000000000000100000000000000000000000000000100; // D (0x0000000100000004) 
//    12'he45 : LOC <=          63'b000000000000000000000000000001000000000000000000000000000000100; // D (0x0000000200000004) 
//    12'hbd4 : LOC <=          63'b000000000000000000000000000010000000000000000000000000000000100; // D (0x0000000400000004) 
//    12'h0f6 : LOC <=          63'b000000000000000000000000000100000000000000000000000000000000100; // D (0x0000000800000004) 
//    12'h38b : LOC <=          63'b000000000000000000000000001000000000000000000000000000000000100; // D (0x0000001000000004) 
//    12'h571 : LOC <=          63'b000000000000000000000000010000000000000000000000000000000000100; // D (0x0000002000000004) 
//    12'h885 : LOC <=          63'b000000000000000000000000100000000000000000000000000000000000100; // D (0x0000004000000004) 
//    12'h654 : LOC <=          63'b000000000000000000000001000000000000000000000000000000000000100; // D (0x0000008000000004) 
//    12'hecf : LOC <=          63'b000000000000000000000010000000000000000000000000000000000000100; // D (0x0000010000000004) 
//    12'hac0 : LOC <=          63'b000000000000000000000100000000000000000000000000000000000000100; // D (0x0000020000000004) 
//    12'h2de : LOC <=          63'b000000000000000000001000000000000000000000000000000000000000100; // D (0x0000040000000004) 
//    12'h7db : LOC <=          63'b000000000000000000010000000000000000000000000000000000000000100; // D (0x0000080000000004) 
//    12'hdd1 : LOC <=          63'b000000000000000000100000000000000000000000000000000000000000100; // D (0x0000100000000004) 
//    12'hcfc : LOC <=          63'b000000000000000001000000000000000000000000000000000000000000100; // D (0x0000200000000004) 
//    12'hea6 : LOC <=          63'b000000000000000010000000000000000000000000000000000000000000100; // D (0x0000400000000004) 
//    12'ha12 : LOC <=          63'b000000000000000100000000000000000000000000000000000000000000100; // D (0x0000800000000004) 
//    12'h37a : LOC <=          63'b000000000000001000000000000000000000000000000000000000000000100; // D (0x0001000000000004) 
//    12'h493 : LOC <=          63'b000000000000010000000000000000000000000000000000000000000000100; // D (0x0002000000000004) 
//    12'hb41 : LOC <=          63'b000000000000100000000000000000000000000000000000000000000000100; // D (0x0004000000000004) 
//    12'h1dc : LOC <=          63'b000000000001000000000000000000000000000000000000000000000000100; // D (0x0008000000000004) 
//    12'h1df : LOC <=          63'b000000000010000000000000000000000000000000000000000000000000100; // D (0x0010000000000004) 
//    12'h1d9 : LOC <=          63'b000000000100000000000000000000000000000000000000000000000000100; // D (0x0020000000000004) 
//    12'h1d5 : LOC <=          63'b000000001000000000000000000000000000000000000000000000000000100; // D (0x0040000000000004) 
//    12'h1cd : LOC <=          63'b000000010000000000000000000000000000000000000000000000000000100; // D (0x0080000000000004) 
//    12'h1fd : LOC <=          63'b000000100000000000000000000000000000000000000000000000000000100; // D (0x0100000000000004) 
//    12'h19d : LOC <=          63'b000001000000000000000000000000000000000000000000000000000000100; // D (0x0200000000000004) 
//    12'h15d : LOC <=          63'b000010000000000000000000000000000000000000000000000000000000100; // D (0x0400000000000004) 
//    12'h0dd : LOC <=          63'b000100000000000000000000000000000000000000000000000000000000100; // D (0x0800000000000004) 
//    12'h3dd : LOC <=          63'b001000000000000000000000000000000000000000000000000000000000100; // D (0x1000000000000004) 
//    12'h5dd : LOC <=          63'b010000000000000000000000000000000000000000000000000000000000100; // D (0x2000000000000004) 
//    12'h9dd : LOC <=          63'b100000000000000000000000000000000000000000000000000000000000100; // D (0x4000000000000004) 
    12'h683 : LOC <=          63'b000000000000000000000000000000000000000000000000000000000001001; // D (0x0000000000000009) 
    12'h9c8 : LOC <=          63'b000000000000000000000000000000000000000000000000000000000001010; // D (0x000000000000000a) 
    12'h267 : LOC <=          63'b000000000000000000000000000000000000000000000000000000000001100; // D (0x000000000000000c) 
    12'h3ba : LOC <=          63'b000000000000000000000000000000000000000000000000000000000001000; // S (0x0000000000000008) 
//    12'h4ce : LOC <=          63'b000000000000000000000000000000000000000000000000000000000011000; // D (0x0000000000000018) 
//    12'hd52 : LOC <=          63'b000000000000000000000000000000000000000000000000000000000101000; // D (0x0000000000000028) 
//    12'hb53 : LOC <=          63'b000000000000000000000000000000000000000000000000000000001001000; // D (0x0000000000000048) 
//    12'h751 : LOC <=          63'b000000000000000000000000000000000000000000000000000000010001000; // D (0x0000000000000088) 
//    12'ha6c : LOC <=          63'b000000000000000000000000000000000000000000000000000000100001000; // D (0x0000000000000108) 
//    12'h52f : LOC <=          63'b000000000000000000000000000000000000000000000000000001000001000; // D (0x0000000000000208) 
//    12'he90 : LOC <=          63'b000000000000000000000000000000000000000000000000000010000001000; // D (0x0000000000000408) 
//    12'hcd7 : LOC <=          63'b000000000000000000000000000000000000000000000000000100000001000; // D (0x0000000000000808) 
//    12'h859 : LOC <=          63'b000000000000000000000000000000000000000000000000001000000001000; // D (0x0000000000001008) 
//    12'h145 : LOC <=          63'b000000000000000000000000000000000000000000000000010000000001000; // D (0x0000000000002008) 
//    12'h644 : LOC <=          63'b000000000000000000000000000000000000000000000000100000000001000; // D (0x0000000000004008) 
//    12'h846 : LOC <=          63'b000000000000000000000000000000000000000000000001000000000001000; // D (0x0000000000008008) 
//    12'h17b : LOC <=          63'b000000000000000000000000000000000000000000000010000000000001000; // D (0x0000000000010008) 
//    12'h638 : LOC <=          63'b000000000000000000000000000000000000000000000100000000000001000; // D (0x0000000000020008) 
//    12'h8be : LOC <=          63'b000000000000000000000000000000000000000000001000000000000001000; // D (0x0000000000040008) 
//    12'h08b : LOC <=          63'b000000000000000000000000000000000000000000010000000000000001000; // D (0x0000000000080008) 
//    12'h5d8 : LOC <=          63'b000000000000000000000000000000000000000000100000000000000001000; // D (0x0000000000100008) 
//    12'hf7e : LOC <=          63'b000000000000000000000000000000000000000001000000000000000001000; // D (0x0000000000200008) 
//    12'hf0b : LOC <=          63'b000000000000000000000000000000000000000010000000000000000001000; // D (0x0000000000400008) 
//    12'hfe1 : LOC <=          63'b000000000000000000000000000000000000000100000000000000000001000; // D (0x0000000000800008) 
//    12'he35 : LOC <=          63'b000000000000000000000000000000000000001000000000000000000001000; // D (0x0000000001000008) 
//    12'hd9d : LOC <=          63'b000000000000000000000000000000000000010000000000000000000001000; // D (0x0000000002000008) 
//    12'hacd : LOC <=          63'b000000000000000000000000000000000000100000000000000000000001000; // D (0x0000000004000008) 
//    12'h46d : LOC <=          63'b000000000000000000000000000000000001000000000000000000000001000; // D (0x0000000008000008) 
//    12'hc14 : LOC <=          63'b000000000000000000000000000000000010000000000000000000000001000; // D (0x0000000010000008) 
//    12'h9df : LOC <=          63'b000000000000000000000000000000000100000000000000000000000001000; // D (0x0000000020000008) 
//    12'h249 : LOC <=          63'b000000000000000000000000000000001000000000000000000000000001000; // D (0x0000000040000008) 
//    12'h05c : LOC <=          63'b000000000000000000000000000000010000000000000000000000000001000; // D (0x0000000080000008) 
//    12'h476 : LOC <=          63'b000000000000000000000000000000100000000000000000000000000001000; // D (0x0000000100000008) 
//    12'hc22 : LOC <=          63'b000000000000000000000000000001000000000000000000000000000001000; // D (0x0000000200000008) 
//    12'h9b3 : LOC <=          63'b000000000000000000000000000010000000000000000000000000000001000; // D (0x0000000400000008) 
//    12'h291 : LOC <=          63'b000000000000000000000000000100000000000000000000000000000001000; // D (0x0000000800000008) 
//    12'h1ec : LOC <=          63'b000000000000000000000000001000000000000000000000000000000001000; // D (0x0000001000000008) 
//    12'h716 : LOC <=          63'b000000000000000000000000010000000000000000000000000000000001000; // D (0x0000002000000008) 
//    12'hae2 : LOC <=          63'b000000000000000000000000100000000000000000000000000000000001000; // D (0x0000004000000008) 
//    12'h433 : LOC <=          63'b000000000000000000000001000000000000000000000000000000000001000; // D (0x0000008000000008) 
//    12'hca8 : LOC <=          63'b000000000000000000000010000000000000000000000000000000000001000; // D (0x0000010000000008) 
//    12'h8a7 : LOC <=          63'b000000000000000000000100000000000000000000000000000000000001000; // D (0x0000020000000008) 
//    12'h0b9 : LOC <=          63'b000000000000000000001000000000000000000000000000000000000001000; // D (0x0000040000000008) 
//    12'h5bc : LOC <=          63'b000000000000000000010000000000000000000000000000000000000001000; // D (0x0000080000000008) 
//    12'hfb6 : LOC <=          63'b000000000000000000100000000000000000000000000000000000000001000; // D (0x0000100000000008) 
//    12'he9b : LOC <=          63'b000000000000000001000000000000000000000000000000000000000001000; // D (0x0000200000000008) 
//    12'hcc1 : LOC <=          63'b000000000000000010000000000000000000000000000000000000000001000; // D (0x0000400000000008) 
//    12'h875 : LOC <=          63'b000000000000000100000000000000000000000000000000000000000001000; // D (0x0000800000000008) 
//    12'h11d : LOC <=          63'b000000000000001000000000000000000000000000000000000000000001000; // D (0x0001000000000008) 
//    12'h6f4 : LOC <=          63'b000000000000010000000000000000000000000000000000000000000001000; // D (0x0002000000000008) 
//    12'h926 : LOC <=          63'b000000000000100000000000000000000000000000000000000000000001000; // D (0x0004000000000008) 
//    12'h3bb : LOC <=          63'b000000000001000000000000000000000000000000000000000000000001000; // D (0x0008000000000008) 
//    12'h3b8 : LOC <=          63'b000000000010000000000000000000000000000000000000000000000001000; // D (0x0010000000000008) 
//    12'h3be : LOC <=          63'b000000000100000000000000000000000000000000000000000000000001000; // D (0x0020000000000008) 
//    12'h3b2 : LOC <=          63'b000000001000000000000000000000000000000000000000000000000001000; // D (0x0040000000000008) 
//    12'h3aa : LOC <=          63'b000000010000000000000000000000000000000000000000000000000001000; // D (0x0080000000000008) 
//    12'h39a : LOC <=          63'b000000100000000000000000000000000000000000000000000000000001000; // D (0x0100000000000008) 
//    12'h3fa : LOC <=          63'b000001000000000000000000000000000000000000000000000000000001000; // D (0x0200000000000008) 
//    12'h33a : LOC <=          63'b000010000000000000000000000000000000000000000000000000000001000; // D (0x0400000000000008) 
//    12'h2ba : LOC <=          63'b000100000000000000000000000000000000000000000000000000000001000; // D (0x0800000000000008) 
//    12'h1ba : LOC <=          63'b001000000000000000000000000000000000000000000000000000000001000; // D (0x1000000000000008) 
//    12'h7ba : LOC <=          63'b010000000000000000000000000000000000000000000000000000000001000; // D (0x2000000000000008) 
//    12'hbba : LOC <=          63'b100000000000000000000000000000000000000000000000000000000001000; // D (0x4000000000000008) 
    12'h24d : LOC <=          63'b000000000000000000000000000000000000000000000000000000000010001; // D (0x0000000000000011) 
    12'hd06 : LOC <=          63'b000000000000000000000000000000000000000000000000000000000010010; // D (0x0000000000000012) 
    12'h6a9 : LOC <=          63'b000000000000000000000000000000000000000000000000000000000010100; // D (0x0000000000000014) 
    12'h4ce : LOC <=          63'b000000000000000000000000000000000000000000000000000000000011000; // D (0x0000000000000018) 
    12'h774 : LOC <=          63'b000000000000000000000000000000000000000000000000000000000010000; // S (0x0000000000000010) 
//    12'h99c : LOC <=          63'b000000000000000000000000000000000000000000000000000000000110000; // D (0x0000000000000030) 
//    12'hf9d : LOC <=          63'b000000000000000000000000000000000000000000000000000000001010000; // D (0x0000000000000050) 
//    12'h39f : LOC <=          63'b000000000000000000000000000000000000000000000000000000010010000; // D (0x0000000000000090) 
//    12'hea2 : LOC <=          63'b000000000000000000000000000000000000000000000000000000100010000; // D (0x0000000000000110) 
//    12'h1e1 : LOC <=          63'b000000000000000000000000000000000000000000000000000001000010000; // D (0x0000000000000210) 
//    12'ha5e : LOC <=          63'b000000000000000000000000000000000000000000000000000010000010000; // D (0x0000000000000410) 
//    12'h819 : LOC <=          63'b000000000000000000000000000000000000000000000000000100000010000; // D (0x0000000000000810) 
//    12'hc97 : LOC <=          63'b000000000000000000000000000000000000000000000000001000000010000; // D (0x0000000000001010) 
//    12'h58b : LOC <=          63'b000000000000000000000000000000000000000000000000010000000010000; // D (0x0000000000002010) 
//    12'h28a : LOC <=          63'b000000000000000000000000000000000000000000000000100000000010000; // D (0x0000000000004010) 
//    12'hc88 : LOC <=          63'b000000000000000000000000000000000000000000000001000000000010000; // D (0x0000000000008010) 
//    12'h5b5 : LOC <=          63'b000000000000000000000000000000000000000000000010000000000010000; // D (0x0000000000010010) 
//    12'h2f6 : LOC <=          63'b000000000000000000000000000000000000000000000100000000000010000; // D (0x0000000000020010) 
//    12'hc70 : LOC <=          63'b000000000000000000000000000000000000000000001000000000000010000; // D (0x0000000000040010) 
//    12'h445 : LOC <=          63'b000000000000000000000000000000000000000000010000000000000010000; // D (0x0000000000080010) 
//    12'h116 : LOC <=          63'b000000000000000000000000000000000000000000100000000000000010000; // D (0x0000000000100010) 
//    12'hbb0 : LOC <=          63'b000000000000000000000000000000000000000001000000000000000010000; // D (0x0000000000200010) 
//    12'hbc5 : LOC <=          63'b000000000000000000000000000000000000000010000000000000000010000; // D (0x0000000000400010) 
//    12'hb2f : LOC <=          63'b000000000000000000000000000000000000000100000000000000000010000; // D (0x0000000000800010) 
//    12'hafb : LOC <=          63'b000000000000000000000000000000000000001000000000000000000010000; // D (0x0000000001000010) 
//    12'h953 : LOC <=          63'b000000000000000000000000000000000000010000000000000000000010000; // D (0x0000000002000010) 
//    12'he03 : LOC <=          63'b000000000000000000000000000000000000100000000000000000000010000; // D (0x0000000004000010) 
//    12'h0a3 : LOC <=          63'b000000000000000000000000000000000001000000000000000000000010000; // D (0x0000000008000010) 
//    12'h8da : LOC <=          63'b000000000000000000000000000000000010000000000000000000000010000; // D (0x0000000010000010) 
//    12'hd11 : LOC <=          63'b000000000000000000000000000000000100000000000000000000000010000; // D (0x0000000020000010) 
//    12'h687 : LOC <=          63'b000000000000000000000000000000001000000000000000000000000010000; // D (0x0000000040000010) 
//    12'h492 : LOC <=          63'b000000000000000000000000000000010000000000000000000000000010000; // D (0x0000000080000010) 
//    12'h0b8 : LOC <=          63'b000000000000000000000000000000100000000000000000000000000010000; // D (0x0000000100000010) 
//    12'h8ec : LOC <=          63'b000000000000000000000000000001000000000000000000000000000010000; // D (0x0000000200000010) 
//    12'hd7d : LOC <=          63'b000000000000000000000000000010000000000000000000000000000010000; // D (0x0000000400000010) 
//    12'h65f : LOC <=          63'b000000000000000000000000000100000000000000000000000000000010000; // D (0x0000000800000010) 
//    12'h522 : LOC <=          63'b000000000000000000000000001000000000000000000000000000000010000; // D (0x0000001000000010) 
//    12'h3d8 : LOC <=          63'b000000000000000000000000010000000000000000000000000000000010000; // D (0x0000002000000010) 
//    12'he2c : LOC <=          63'b000000000000000000000000100000000000000000000000000000000010000; // D (0x0000004000000010) 
//    12'h0fd : LOC <=          63'b000000000000000000000001000000000000000000000000000000000010000; // D (0x0000008000000010) 
//    12'h866 : LOC <=          63'b000000000000000000000010000000000000000000000000000000000010000; // D (0x0000010000000010) 
//    12'hc69 : LOC <=          63'b000000000000000000000100000000000000000000000000000000000010000; // D (0x0000020000000010) 
//    12'h477 : LOC <=          63'b000000000000000000001000000000000000000000000000000000000010000; // D (0x0000040000000010) 
//    12'h172 : LOC <=          63'b000000000000000000010000000000000000000000000000000000000010000; // D (0x0000080000000010) 
//    12'hb78 : LOC <=          63'b000000000000000000100000000000000000000000000000000000000010000; // D (0x0000100000000010) 
//    12'ha55 : LOC <=          63'b000000000000000001000000000000000000000000000000000000000010000; // D (0x0000200000000010) 
//    12'h80f : LOC <=          63'b000000000000000010000000000000000000000000000000000000000010000; // D (0x0000400000000010) 
//    12'hcbb : LOC <=          63'b000000000000000100000000000000000000000000000000000000000010000; // D (0x0000800000000010) 
//    12'h5d3 : LOC <=          63'b000000000000001000000000000000000000000000000000000000000010000; // D (0x0001000000000010) 
//    12'h23a : LOC <=          63'b000000000000010000000000000000000000000000000000000000000010000; // D (0x0002000000000010) 
//    12'hde8 : LOC <=          63'b000000000000100000000000000000000000000000000000000000000010000; // D (0x0004000000000010) 
//    12'h775 : LOC <=          63'b000000000001000000000000000000000000000000000000000000000010000; // D (0x0008000000000010) 
//    12'h776 : LOC <=          63'b000000000010000000000000000000000000000000000000000000000010000; // D (0x0010000000000010) 
//    12'h770 : LOC <=          63'b000000000100000000000000000000000000000000000000000000000010000; // D (0x0020000000000010) 
//    12'h77c : LOC <=          63'b000000001000000000000000000000000000000000000000000000000010000; // D (0x0040000000000010) 
//    12'h764 : LOC <=          63'b000000010000000000000000000000000000000000000000000000000010000; // D (0x0080000000000010) 
//    12'h754 : LOC <=          63'b000000100000000000000000000000000000000000000000000000000010000; // D (0x0100000000000010) 
//    12'h734 : LOC <=          63'b000001000000000000000000000000000000000000000000000000000010000; // D (0x0200000000000010) 
//    12'h7f4 : LOC <=          63'b000010000000000000000000000000000000000000000000000000000010000; // D (0x0400000000000010) 
//    12'h674 : LOC <=          63'b000100000000000000000000000000000000000000000000000000000010000; // D (0x0800000000000010) 
//    12'h574 : LOC <=          63'b001000000000000000000000000000000000000000000000000000000010000; // D (0x1000000000000010) 
//    12'h374 : LOC <=          63'b010000000000000000000000000000000000000000000000000000000010000; // D (0x2000000000000010) 
//    12'hf74 : LOC <=          63'b100000000000000000000000000000000000000000000000000000000010000; // D (0x4000000000000010) 
    12'hbd1 : LOC <=          63'b000000000000000000000000000000000000000000000000000000000100001; // D (0x0000000000000021) 
    12'h49a : LOC <=          63'b000000000000000000000000000000000000000000000000000000000100010; // D (0x0000000000000022) 
    12'hf35 : LOC <=          63'b000000000000000000000000000000000000000000000000000000000100100; // D (0x0000000000000024) 
    12'hd52 : LOC <=          63'b000000000000000000000000000000000000000000000000000000000101000; // D (0x0000000000000028) 
    12'h99c : LOC <=          63'b000000000000000000000000000000000000000000000000000000000110000; // D (0x0000000000000030) 
    12'hee8 : LOC <=          63'b000000000000000000000000000000000000000000000000000000000100000; // S (0x0000000000000020) 
//    12'h601 : LOC <=          63'b000000000000000000000000000000000000000000000000000000001100000; // D (0x0000000000000060) 
//    12'ha03 : LOC <=          63'b000000000000000000000000000000000000000000000000000000010100000; // D (0x00000000000000a0) 
//    12'h73e : LOC <=          63'b000000000000000000000000000000000000000000000000000000100100000; // D (0x0000000000000120) 
//    12'h87d : LOC <=          63'b000000000000000000000000000000000000000000000000000001000100000; // D (0x0000000000000220) 
//    12'h3c2 : LOC <=          63'b000000000000000000000000000000000000000000000000000010000100000; // D (0x0000000000000420) 
//    12'h185 : LOC <=          63'b000000000000000000000000000000000000000000000000000100000100000; // D (0x0000000000000820) 
//    12'h50b : LOC <=          63'b000000000000000000000000000000000000000000000000001000000100000; // D (0x0000000000001020) 
//    12'hc17 : LOC <=          63'b000000000000000000000000000000000000000000000000010000000100000; // D (0x0000000000002020) 
//    12'hb16 : LOC <=          63'b000000000000000000000000000000000000000000000000100000000100000; // D (0x0000000000004020) 
//    12'h514 : LOC <=          63'b000000000000000000000000000000000000000000000001000000000100000; // D (0x0000000000008020) 
//    12'hc29 : LOC <=          63'b000000000000000000000000000000000000000000000010000000000100000; // D (0x0000000000010020) 
//    12'hb6a : LOC <=          63'b000000000000000000000000000000000000000000000100000000000100000; // D (0x0000000000020020) 
//    12'h5ec : LOC <=          63'b000000000000000000000000000000000000000000001000000000000100000; // D (0x0000000000040020) 
//    12'hdd9 : LOC <=          63'b000000000000000000000000000000000000000000010000000000000100000; // D (0x0000000000080020) 
//    12'h88a : LOC <=          63'b000000000000000000000000000000000000000000100000000000000100000; // D (0x0000000000100020) 
//    12'h22c : LOC <=          63'b000000000000000000000000000000000000000001000000000000000100000; // D (0x0000000000200020) 
//    12'h259 : LOC <=          63'b000000000000000000000000000000000000000010000000000000000100000; // D (0x0000000000400020) 
//    12'h2b3 : LOC <=          63'b000000000000000000000000000000000000000100000000000000000100000; // D (0x0000000000800020) 
//    12'h367 : LOC <=          63'b000000000000000000000000000000000000001000000000000000000100000; // D (0x0000000001000020) 
//    12'h0cf : LOC <=          63'b000000000000000000000000000000000000010000000000000000000100000; // D (0x0000000002000020) 
//    12'h79f : LOC <=          63'b000000000000000000000000000000000000100000000000000000000100000; // D (0x0000000004000020) 
//    12'h93f : LOC <=          63'b000000000000000000000000000000000001000000000000000000000100000; // D (0x0000000008000020) 
//    12'h146 : LOC <=          63'b000000000000000000000000000000000010000000000000000000000100000; // D (0x0000000010000020) 
//    12'h48d : LOC <=          63'b000000000000000000000000000000000100000000000000000000000100000; // D (0x0000000020000020) 
//    12'hf1b : LOC <=          63'b000000000000000000000000000000001000000000000000000000000100000; // D (0x0000000040000020) 
//    12'hd0e : LOC <=          63'b000000000000000000000000000000010000000000000000000000000100000; // D (0x0000000080000020) 
//    12'h924 : LOC <=          63'b000000000000000000000000000000100000000000000000000000000100000; // D (0x0000000100000020) 
//    12'h170 : LOC <=          63'b000000000000000000000000000001000000000000000000000000000100000; // D (0x0000000200000020) 
//    12'h4e1 : LOC <=          63'b000000000000000000000000000010000000000000000000000000000100000; // D (0x0000000400000020) 
//    12'hfc3 : LOC <=          63'b000000000000000000000000000100000000000000000000000000000100000; // D (0x0000000800000020) 
//    12'hcbe : LOC <=          63'b000000000000000000000000001000000000000000000000000000000100000; // D (0x0000001000000020) 
//    12'ha44 : LOC <=          63'b000000000000000000000000010000000000000000000000000000000100000; // D (0x0000002000000020) 
//    12'h7b0 : LOC <=          63'b000000000000000000000000100000000000000000000000000000000100000; // D (0x0000004000000020) 
//    12'h961 : LOC <=          63'b000000000000000000000001000000000000000000000000000000000100000; // D (0x0000008000000020) 
//    12'h1fa : LOC <=          63'b000000000000000000000010000000000000000000000000000000000100000; // D (0x0000010000000020) 
//    12'h5f5 : LOC <=          63'b000000000000000000000100000000000000000000000000000000000100000; // D (0x0000020000000020) 
//    12'hdeb : LOC <=          63'b000000000000000000001000000000000000000000000000000000000100000; // D (0x0000040000000020) 
//    12'h8ee : LOC <=          63'b000000000000000000010000000000000000000000000000000000000100000; // D (0x0000080000000020) 
//    12'h2e4 : LOC <=          63'b000000000000000000100000000000000000000000000000000000000100000; // D (0x0000100000000020) 
//    12'h3c9 : LOC <=          63'b000000000000000001000000000000000000000000000000000000000100000; // D (0x0000200000000020) 
//    12'h193 : LOC <=          63'b000000000000000010000000000000000000000000000000000000000100000; // D (0x0000400000000020) 
//    12'h527 : LOC <=          63'b000000000000000100000000000000000000000000000000000000000100000; // D (0x0000800000000020) 
//    12'hc4f : LOC <=          63'b000000000000001000000000000000000000000000000000000000000100000; // D (0x0001000000000020) 
//    12'hba6 : LOC <=          63'b000000000000010000000000000000000000000000000000000000000100000; // D (0x0002000000000020) 
//    12'h474 : LOC <=          63'b000000000000100000000000000000000000000000000000000000000100000; // D (0x0004000000000020) 
//    12'hee9 : LOC <=          63'b000000000001000000000000000000000000000000000000000000000100000; // D (0x0008000000000020) 
//    12'heea : LOC <=          63'b000000000010000000000000000000000000000000000000000000000100000; // D (0x0010000000000020) 
//    12'heec : LOC <=          63'b000000000100000000000000000000000000000000000000000000000100000; // D (0x0020000000000020) 
//    12'hee0 : LOC <=          63'b000000001000000000000000000000000000000000000000000000000100000; // D (0x0040000000000020) 
//    12'hef8 : LOC <=          63'b000000010000000000000000000000000000000000000000000000000100000; // D (0x0080000000000020) 
//    12'hec8 : LOC <=          63'b000000100000000000000000000000000000000000000000000000000100000; // D (0x0100000000000020) 
//    12'hea8 : LOC <=          63'b000001000000000000000000000000000000000000000000000000000100000; // D (0x0200000000000020) 
//    12'he68 : LOC <=          63'b000010000000000000000000000000000000000000000000000000000100000; // D (0x0400000000000020) 
//    12'hfe8 : LOC <=          63'b000100000000000000000000000000000000000000000000000000000100000; // D (0x0800000000000020) 
//    12'hce8 : LOC <=          63'b001000000000000000000000000000000000000000000000000000000100000; // D (0x1000000000000020) 
//    12'hae8 : LOC <=          63'b010000000000000000000000000000000000000000000000000000000100000; // D (0x2000000000000020) 
//    12'h6e8 : LOC <=          63'b100000000000000000000000000000000000000000000000000000000100000; // D (0x4000000000000020) 
    12'hdd0 : LOC <=          63'b000000000000000000000000000000000000000000000000000000001000001; // D (0x0000000000000041) 
    12'h29b : LOC <=          63'b000000000000000000000000000000000000000000000000000000001000010; // D (0x0000000000000042) 
    12'h934 : LOC <=          63'b000000000000000000000000000000000000000000000000000000001000100; // D (0x0000000000000044) 
    12'hb53 : LOC <=          63'b000000000000000000000000000000000000000000000000000000001001000; // D (0x0000000000000048) 
    12'hf9d : LOC <=          63'b000000000000000000000000000000000000000000000000000000001010000; // D (0x0000000000000050) 
    12'h601 : LOC <=          63'b000000000000000000000000000000000000000000000000000000001100000; // D (0x0000000000000060) 
    12'h8e9 : LOC <=          63'b000000000000000000000000000000000000000000000000000000001000000; // S (0x0000000000000040) 
//    12'hc02 : LOC <=          63'b000000000000000000000000000000000000000000000000000000011000000; // D (0x00000000000000c0) 
//    12'h13f : LOC <=          63'b000000000000000000000000000000000000000000000000000000101000000; // D (0x0000000000000140) 
//    12'he7c : LOC <=          63'b000000000000000000000000000000000000000000000000000001001000000; // D (0x0000000000000240) 
//    12'h5c3 : LOC <=          63'b000000000000000000000000000000000000000000000000000010001000000; // D (0x0000000000000440) 
//    12'h784 : LOC <=          63'b000000000000000000000000000000000000000000000000000100001000000; // D (0x0000000000000840) 
//    12'h30a : LOC <=          63'b000000000000000000000000000000000000000000000000001000001000000; // D (0x0000000000001040) 
//    12'ha16 : LOC <=          63'b000000000000000000000000000000000000000000000000010000001000000; // D (0x0000000000002040) 
//    12'hd17 : LOC <=          63'b000000000000000000000000000000000000000000000000100000001000000; // D (0x0000000000004040) 
//    12'h315 : LOC <=          63'b000000000000000000000000000000000000000000000001000000001000000; // D (0x0000000000008040) 
//    12'ha28 : LOC <=          63'b000000000000000000000000000000000000000000000010000000001000000; // D (0x0000000000010040) 
//    12'hd6b : LOC <=          63'b000000000000000000000000000000000000000000000100000000001000000; // D (0x0000000000020040) 
//    12'h3ed : LOC <=          63'b000000000000000000000000000000000000000000001000000000001000000; // D (0x0000000000040040) 
//    12'hbd8 : LOC <=          63'b000000000000000000000000000000000000000000010000000000001000000; // D (0x0000000000080040) 
//    12'he8b : LOC <=          63'b000000000000000000000000000000000000000000100000000000001000000; // D (0x0000000000100040) 
//    12'h42d : LOC <=          63'b000000000000000000000000000000000000000001000000000000001000000; // D (0x0000000000200040) 
//    12'h458 : LOC <=          63'b000000000000000000000000000000000000000010000000000000001000000; // D (0x0000000000400040) 
//    12'h4b2 : LOC <=          63'b000000000000000000000000000000000000000100000000000000001000000; // D (0x0000000000800040) 
//    12'h566 : LOC <=          63'b000000000000000000000000000000000000001000000000000000001000000; // D (0x0000000001000040) 
//    12'h6ce : LOC <=          63'b000000000000000000000000000000000000010000000000000000001000000; // D (0x0000000002000040) 
//    12'h19e : LOC <=          63'b000000000000000000000000000000000000100000000000000000001000000; // D (0x0000000004000040) 
//    12'hf3e : LOC <=          63'b000000000000000000000000000000000001000000000000000000001000000; // D (0x0000000008000040) 
//    12'h747 : LOC <=          63'b000000000000000000000000000000000010000000000000000000001000000; // D (0x0000000010000040) 
//    12'h28c : LOC <=          63'b000000000000000000000000000000000100000000000000000000001000000; // D (0x0000000020000040) 
//    12'h91a : LOC <=          63'b000000000000000000000000000000001000000000000000000000001000000; // D (0x0000000040000040) 
//    12'hb0f : LOC <=          63'b000000000000000000000000000000010000000000000000000000001000000; // D (0x0000000080000040) 
//    12'hf25 : LOC <=          63'b000000000000000000000000000000100000000000000000000000001000000; // D (0x0000000100000040) 
//    12'h771 : LOC <=          63'b000000000000000000000000000001000000000000000000000000001000000; // D (0x0000000200000040) 
//    12'h2e0 : LOC <=          63'b000000000000000000000000000010000000000000000000000000001000000; // D (0x0000000400000040) 
//    12'h9c2 : LOC <=          63'b000000000000000000000000000100000000000000000000000000001000000; // D (0x0000000800000040) 
//    12'habf : LOC <=          63'b000000000000000000000000001000000000000000000000000000001000000; // D (0x0000001000000040) 
//    12'hc45 : LOC <=          63'b000000000000000000000000010000000000000000000000000000001000000; // D (0x0000002000000040) 
//    12'h1b1 : LOC <=          63'b000000000000000000000000100000000000000000000000000000001000000; // D (0x0000004000000040) 
//    12'hf60 : LOC <=          63'b000000000000000000000001000000000000000000000000000000001000000; // D (0x0000008000000040) 
//    12'h7fb : LOC <=          63'b000000000000000000000010000000000000000000000000000000001000000; // D (0x0000010000000040) 
//    12'h3f4 : LOC <=          63'b000000000000000000000100000000000000000000000000000000001000000; // D (0x0000020000000040) 
//    12'hbea : LOC <=          63'b000000000000000000001000000000000000000000000000000000001000000; // D (0x0000040000000040) 
//    12'heef : LOC <=          63'b000000000000000000010000000000000000000000000000000000001000000; // D (0x0000080000000040) 
//    12'h4e5 : LOC <=          63'b000000000000000000100000000000000000000000000000000000001000000; // D (0x0000100000000040) 
//    12'h5c8 : LOC <=          63'b000000000000000001000000000000000000000000000000000000001000000; // D (0x0000200000000040) 
//    12'h792 : LOC <=          63'b000000000000000010000000000000000000000000000000000000001000000; // D (0x0000400000000040) 
//    12'h326 : LOC <=          63'b000000000000000100000000000000000000000000000000000000001000000; // D (0x0000800000000040) 
//    12'ha4e : LOC <=          63'b000000000000001000000000000000000000000000000000000000001000000; // D (0x0001000000000040) 
//    12'hda7 : LOC <=          63'b000000000000010000000000000000000000000000000000000000001000000; // D (0x0002000000000040) 
//    12'h275 : LOC <=          63'b000000000000100000000000000000000000000000000000000000001000000; // D (0x0004000000000040) 
//    12'h8e8 : LOC <=          63'b000000000001000000000000000000000000000000000000000000001000000; // D (0x0008000000000040) 
//    12'h8eb : LOC <=          63'b000000000010000000000000000000000000000000000000000000001000000; // D (0x0010000000000040) 
//    12'h8ed : LOC <=          63'b000000000100000000000000000000000000000000000000000000001000000; // D (0x0020000000000040) 
//    12'h8e1 : LOC <=          63'b000000001000000000000000000000000000000000000000000000001000000; // D (0x0040000000000040) 
//    12'h8f9 : LOC <=          63'b000000010000000000000000000000000000000000000000000000001000000; // D (0x0080000000000040) 
//    12'h8c9 : LOC <=          63'b000000100000000000000000000000000000000000000000000000001000000; // D (0x0100000000000040) 
//    12'h8a9 : LOC <=          63'b000001000000000000000000000000000000000000000000000000001000000; // D (0x0200000000000040) 
//    12'h869 : LOC <=          63'b000010000000000000000000000000000000000000000000000000001000000; // D (0x0400000000000040) 
//    12'h9e9 : LOC <=          63'b000100000000000000000000000000000000000000000000000000001000000; // D (0x0800000000000040) 
//    12'hae9 : LOC <=          63'b001000000000000000000000000000000000000000000000000000001000000; // D (0x1000000000000040) 
//    12'hce9 : LOC <=          63'b010000000000000000000000000000000000000000000000000000001000000; // D (0x2000000000000040) 
//    12'h0e9 : LOC <=          63'b100000000000000000000000000000000000000000000000000000001000000; // D (0x4000000000000040) 
    12'h1d2 : LOC <=          63'b000000000000000000000000000000000000000000000000000000010000001; // D (0x0000000000000081) 
    12'he99 : LOC <=          63'b000000000000000000000000000000000000000000000000000000010000010; // D (0x0000000000000082) 
    12'h536 : LOC <=          63'b000000000000000000000000000000000000000000000000000000010000100; // D (0x0000000000000084) 
    12'h751 : LOC <=          63'b000000000000000000000000000000000000000000000000000000010001000; // D (0x0000000000000088) 
    12'h39f : LOC <=          63'b000000000000000000000000000000000000000000000000000000010010000; // D (0x0000000000000090) 
    12'ha03 : LOC <=          63'b000000000000000000000000000000000000000000000000000000010100000; // D (0x00000000000000a0) 
    12'hc02 : LOC <=          63'b000000000000000000000000000000000000000000000000000000011000000; // D (0x00000000000000c0) 
    12'h4eb : LOC <=          63'b000000000000000000000000000000000000000000000000000000010000000; // S (0x0000000000000080) 
//    12'hd3d : LOC <=          63'b000000000000000000000000000000000000000000000000000000110000000; // D (0x0000000000000180) 
//    12'h27e : LOC <=          63'b000000000000000000000000000000000000000000000000000001010000000; // D (0x0000000000000280) 
//    12'h9c1 : LOC <=          63'b000000000000000000000000000000000000000000000000000010010000000; // D (0x0000000000000480) 
//    12'hb86 : LOC <=          63'b000000000000000000000000000000000000000000000000000100010000000; // D (0x0000000000000880) 
//    12'hf08 : LOC <=          63'b000000000000000000000000000000000000000000000000001000010000000; // D (0x0000000000001080) 
//    12'h614 : LOC <=          63'b000000000000000000000000000000000000000000000000010000010000000; // D (0x0000000000002080) 
//    12'h115 : LOC <=          63'b000000000000000000000000000000000000000000000000100000010000000; // D (0x0000000000004080) 
//    12'hf17 : LOC <=          63'b000000000000000000000000000000000000000000000001000000010000000; // D (0x0000000000008080) 
//    12'h62a : LOC <=          63'b000000000000000000000000000000000000000000000010000000010000000; // D (0x0000000000010080) 
//    12'h169 : LOC <=          63'b000000000000000000000000000000000000000000000100000000010000000; // D (0x0000000000020080) 
//    12'hfef : LOC <=          63'b000000000000000000000000000000000000000000001000000000010000000; // D (0x0000000000040080) 
//    12'h7da : LOC <=          63'b000000000000000000000000000000000000000000010000000000010000000; // D (0x0000000000080080) 
//    12'h289 : LOC <=          63'b000000000000000000000000000000000000000000100000000000010000000; // D (0x0000000000100080) 
//    12'h82f : LOC <=          63'b000000000000000000000000000000000000000001000000000000010000000; // D (0x0000000000200080) 
//    12'h85a : LOC <=          63'b000000000000000000000000000000000000000010000000000000010000000; // D (0x0000000000400080) 
//    12'h8b0 : LOC <=          63'b000000000000000000000000000000000000000100000000000000010000000; // D (0x0000000000800080) 
//    12'h964 : LOC <=          63'b000000000000000000000000000000000000001000000000000000010000000; // D (0x0000000001000080) 
//    12'hacc : LOC <=          63'b000000000000000000000000000000000000010000000000000000010000000; // D (0x0000000002000080) 
//    12'hd9c : LOC <=          63'b000000000000000000000000000000000000100000000000000000010000000; // D (0x0000000004000080) 
//    12'h33c : LOC <=          63'b000000000000000000000000000000000001000000000000000000010000000; // D (0x0000000008000080) 
//    12'hb45 : LOC <=          63'b000000000000000000000000000000000010000000000000000000010000000; // D (0x0000000010000080) 
//    12'he8e : LOC <=          63'b000000000000000000000000000000000100000000000000000000010000000; // D (0x0000000020000080) 
//    12'h518 : LOC <=          63'b000000000000000000000000000000001000000000000000000000010000000; // D (0x0000000040000080) 
//    12'h70d : LOC <=          63'b000000000000000000000000000000010000000000000000000000010000000; // D (0x0000000080000080) 
//    12'h327 : LOC <=          63'b000000000000000000000000000000100000000000000000000000010000000; // D (0x0000000100000080) 
//    12'hb73 : LOC <=          63'b000000000000000000000000000001000000000000000000000000010000000; // D (0x0000000200000080) 
//    12'hee2 : LOC <=          63'b000000000000000000000000000010000000000000000000000000010000000; // D (0x0000000400000080) 
//    12'h5c0 : LOC <=          63'b000000000000000000000000000100000000000000000000000000010000000; // D (0x0000000800000080) 
//    12'h6bd : LOC <=          63'b000000000000000000000000001000000000000000000000000000010000000; // D (0x0000001000000080) 
//    12'h047 : LOC <=          63'b000000000000000000000000010000000000000000000000000000010000000; // D (0x0000002000000080) 
//    12'hdb3 : LOC <=          63'b000000000000000000000000100000000000000000000000000000010000000; // D (0x0000004000000080) 
//    12'h362 : LOC <=          63'b000000000000000000000001000000000000000000000000000000010000000; // D (0x0000008000000080) 
//    12'hbf9 : LOC <=          63'b000000000000000000000010000000000000000000000000000000010000000; // D (0x0000010000000080) 
//    12'hff6 : LOC <=          63'b000000000000000000000100000000000000000000000000000000010000000; // D (0x0000020000000080) 
//    12'h7e8 : LOC <=          63'b000000000000000000001000000000000000000000000000000000010000000; // D (0x0000040000000080) 
//    12'h2ed : LOC <=          63'b000000000000000000010000000000000000000000000000000000010000000; // D (0x0000080000000080) 
//    12'h8e7 : LOC <=          63'b000000000000000000100000000000000000000000000000000000010000000; // D (0x0000100000000080) 
//    12'h9ca : LOC <=          63'b000000000000000001000000000000000000000000000000000000010000000; // D (0x0000200000000080) 
//    12'hb90 : LOC <=          63'b000000000000000010000000000000000000000000000000000000010000000; // D (0x0000400000000080) 
//    12'hf24 : LOC <=          63'b000000000000000100000000000000000000000000000000000000010000000; // D (0x0000800000000080) 
//    12'h64c : LOC <=          63'b000000000000001000000000000000000000000000000000000000010000000; // D (0x0001000000000080) 
//    12'h1a5 : LOC <=          63'b000000000000010000000000000000000000000000000000000000010000000; // D (0x0002000000000080) 
//    12'he77 : LOC <=          63'b000000000000100000000000000000000000000000000000000000010000000; // D (0x0004000000000080) 
//    12'h4ea : LOC <=          63'b000000000001000000000000000000000000000000000000000000010000000; // D (0x0008000000000080) 
//    12'h4e9 : LOC <=          63'b000000000010000000000000000000000000000000000000000000010000000; // D (0x0010000000000080) 
//    12'h4ef : LOC <=          63'b000000000100000000000000000000000000000000000000000000010000000; // D (0x0020000000000080) 
//    12'h4e3 : LOC <=          63'b000000001000000000000000000000000000000000000000000000010000000; // D (0x0040000000000080) 
//    12'h4fb : LOC <=          63'b000000010000000000000000000000000000000000000000000000010000000; // D (0x0080000000000080) 
//    12'h4cb : LOC <=          63'b000000100000000000000000000000000000000000000000000000010000000; // D (0x0100000000000080) 
//    12'h4ab : LOC <=          63'b000001000000000000000000000000000000000000000000000000010000000; // D (0x0200000000000080) 
//    12'h46b : LOC <=          63'b000010000000000000000000000000000000000000000000000000010000000; // D (0x0400000000000080) 
//    12'h5eb : LOC <=          63'b000100000000000000000000000000000000000000000000000000010000000; // D (0x0800000000000080) 
//    12'h6eb : LOC <=          63'b001000000000000000000000000000000000000000000000000000010000000; // D (0x1000000000000080) 
//    12'h0eb : LOC <=          63'b010000000000000000000000000000000000000000000000000000010000000; // D (0x2000000000000080) 
//    12'hceb : LOC <=          63'b100000000000000000000000000000000000000000000000000000010000000; // D (0x4000000000000080) 
    12'hcef : LOC <=          63'b000000000000000000000000000000000000000000000000000000100000001; // D (0x0000000000000101) 
    12'h3a4 : LOC <=          63'b000000000000000000000000000000000000000000000000000000100000010; // D (0x0000000000000102) 
    12'h80b : LOC <=          63'b000000000000000000000000000000000000000000000000000000100000100; // D (0x0000000000000104) 
    12'ha6c : LOC <=          63'b000000000000000000000000000000000000000000000000000000100001000; // D (0x0000000000000108) 
    12'hea2 : LOC <=          63'b000000000000000000000000000000000000000000000000000000100010000; // D (0x0000000000000110) 
    12'h73e : LOC <=          63'b000000000000000000000000000000000000000000000000000000100100000; // D (0x0000000000000120) 
    12'h13f : LOC <=          63'b000000000000000000000000000000000000000000000000000000101000000; // D (0x0000000000000140) 
    12'hd3d : LOC <=          63'b000000000000000000000000000000000000000000000000000000110000000; // D (0x0000000000000180) 
    12'h9d6 : LOC <=          63'b000000000000000000000000000000000000000000000000000000100000000; // S (0x0000000000000100) 
//    12'hf43 : LOC <=          63'b000000000000000000000000000000000000000000000000000001100000000; // D (0x0000000000000300) 
//    12'h4fc : LOC <=          63'b000000000000000000000000000000000000000000000000000010100000000; // D (0x0000000000000500) 
//    12'h6bb : LOC <=          63'b000000000000000000000000000000000000000000000000000100100000000; // D (0x0000000000000900) 
//    12'h235 : LOC <=          63'b000000000000000000000000000000000000000000000000001000100000000; // D (0x0000000000001100) 
//    12'hb29 : LOC <=          63'b000000000000000000000000000000000000000000000000010000100000000; // D (0x0000000000002100) 
//    12'hc28 : LOC <=          63'b000000000000000000000000000000000000000000000000100000100000000; // D (0x0000000000004100) 
//    12'h22a : LOC <=          63'b000000000000000000000000000000000000000000000001000000100000000; // D (0x0000000000008100) 
//    12'hb17 : LOC <=          63'b000000000000000000000000000000000000000000000010000000100000000; // D (0x0000000000010100) 
//    12'hc54 : LOC <=          63'b000000000000000000000000000000000000000000000100000000100000000; // D (0x0000000000020100) 
//    12'h2d2 : LOC <=          63'b000000000000000000000000000000000000000000001000000000100000000; // D (0x0000000000040100) 
//    12'hae7 : LOC <=          63'b000000000000000000000000000000000000000000010000000000100000000; // D (0x0000000000080100) 
//    12'hfb4 : LOC <=          63'b000000000000000000000000000000000000000000100000000000100000000; // D (0x0000000000100100) 
//    12'h512 : LOC <=          63'b000000000000000000000000000000000000000001000000000000100000000; // D (0x0000000000200100) 
//    12'h567 : LOC <=          63'b000000000000000000000000000000000000000010000000000000100000000; // D (0x0000000000400100) 
//    12'h58d : LOC <=          63'b000000000000000000000000000000000000000100000000000000100000000; // D (0x0000000000800100) 
//    12'h459 : LOC <=          63'b000000000000000000000000000000000000001000000000000000100000000; // D (0x0000000001000100) 
//    12'h7f1 : LOC <=          63'b000000000000000000000000000000000000010000000000000000100000000; // D (0x0000000002000100) 
//    12'h0a1 : LOC <=          63'b000000000000000000000000000000000000100000000000000000100000000; // D (0x0000000004000100) 
//    12'he01 : LOC <=          63'b000000000000000000000000000000000001000000000000000000100000000; // D (0x0000000008000100) 
//    12'h678 : LOC <=          63'b000000000000000000000000000000000010000000000000000000100000000; // D (0x0000000010000100) 
//    12'h3b3 : LOC <=          63'b000000000000000000000000000000000100000000000000000000100000000; // D (0x0000000020000100) 
//    12'h825 : LOC <=          63'b000000000000000000000000000000001000000000000000000000100000000; // D (0x0000000040000100) 
//    12'ha30 : LOC <=          63'b000000000000000000000000000000010000000000000000000000100000000; // D (0x0000000080000100) 
//    12'he1a : LOC <=          63'b000000000000000000000000000000100000000000000000000000100000000; // D (0x0000000100000100) 
//    12'h64e : LOC <=          63'b000000000000000000000000000001000000000000000000000000100000000; // D (0x0000000200000100) 
//    12'h3df : LOC <=          63'b000000000000000000000000000010000000000000000000000000100000000; // D (0x0000000400000100) 
//    12'h8fd : LOC <=          63'b000000000000000000000000000100000000000000000000000000100000000; // D (0x0000000800000100) 
//    12'hb80 : LOC <=          63'b000000000000000000000000001000000000000000000000000000100000000; // D (0x0000001000000100) 
//    12'hd7a : LOC <=          63'b000000000000000000000000010000000000000000000000000000100000000; // D (0x0000002000000100) 
//    12'h08e : LOC <=          63'b000000000000000000000000100000000000000000000000000000100000000; // D (0x0000004000000100) 
//    12'he5f : LOC <=          63'b000000000000000000000001000000000000000000000000000000100000000; // D (0x0000008000000100) 
//    12'h6c4 : LOC <=          63'b000000000000000000000010000000000000000000000000000000100000000; // D (0x0000010000000100) 
//    12'h2cb : LOC <=          63'b000000000000000000000100000000000000000000000000000000100000000; // D (0x0000020000000100) 
//    12'had5 : LOC <=          63'b000000000000000000001000000000000000000000000000000000100000000; // D (0x0000040000000100) 
//    12'hfd0 : LOC <=          63'b000000000000000000010000000000000000000000000000000000100000000; // D (0x0000080000000100) 
//    12'h5da : LOC <=          63'b000000000000000000100000000000000000000000000000000000100000000; // D (0x0000100000000100) 
//    12'h4f7 : LOC <=          63'b000000000000000001000000000000000000000000000000000000100000000; // D (0x0000200000000100) 
//    12'h6ad : LOC <=          63'b000000000000000010000000000000000000000000000000000000100000000; // D (0x0000400000000100) 
//    12'h219 : LOC <=          63'b000000000000000100000000000000000000000000000000000000100000000; // D (0x0000800000000100) 
//    12'hb71 : LOC <=          63'b000000000000001000000000000000000000000000000000000000100000000; // D (0x0001000000000100) 
//    12'hc98 : LOC <=          63'b000000000000010000000000000000000000000000000000000000100000000; // D (0x0002000000000100) 
//    12'h34a : LOC <=          63'b000000000000100000000000000000000000000000000000000000100000000; // D (0x0004000000000100) 
//    12'h9d7 : LOC <=          63'b000000000001000000000000000000000000000000000000000000100000000; // D (0x0008000000000100) 
//    12'h9d4 : LOC <=          63'b000000000010000000000000000000000000000000000000000000100000000; // D (0x0010000000000100) 
//    12'h9d2 : LOC <=          63'b000000000100000000000000000000000000000000000000000000100000000; // D (0x0020000000000100) 
//    12'h9de : LOC <=          63'b000000001000000000000000000000000000000000000000000000100000000; // D (0x0040000000000100) 
//    12'h9c6 : LOC <=          63'b000000010000000000000000000000000000000000000000000000100000000; // D (0x0080000000000100) 
//    12'h9f6 : LOC <=          63'b000000100000000000000000000000000000000000000000000000100000000; // D (0x0100000000000100) 
//    12'h996 : LOC <=          63'b000001000000000000000000000000000000000000000000000000100000000; // D (0x0200000000000100) 
//    12'h956 : LOC <=          63'b000010000000000000000000000000000000000000000000000000100000000; // D (0x0400000000000100) 
//    12'h8d6 : LOC <=          63'b000100000000000000000000000000000000000000000000000000100000000; // D (0x0800000000000100) 
//    12'hbd6 : LOC <=          63'b001000000000000000000000000000000000000000000000000000100000000; // D (0x1000000000000100) 
//    12'hdd6 : LOC <=          63'b010000000000000000000000000000000000000000000000000000100000000; // D (0x2000000000000100) 
//    12'h1d6 : LOC <=          63'b100000000000000000000000000000000000000000000000000000100000000; // D (0x4000000000000100) 
    12'h3ac : LOC <=          63'b000000000000000000000000000000000000000000000000000001000000001; // D (0x0000000000000201) 
    12'hce7 : LOC <=          63'b000000000000000000000000000000000000000000000000000001000000010; // D (0x0000000000000202) 
    12'h748 : LOC <=          63'b000000000000000000000000000000000000000000000000000001000000100; // D (0x0000000000000204) 
    12'h52f : LOC <=          63'b000000000000000000000000000000000000000000000000000001000001000; // D (0x0000000000000208) 
    12'h1e1 : LOC <=          63'b000000000000000000000000000000000000000000000000000001000010000; // D (0x0000000000000210) 
    12'h87d : LOC <=          63'b000000000000000000000000000000000000000000000000000001000100000; // D (0x0000000000000220) 
    12'he7c : LOC <=          63'b000000000000000000000000000000000000000000000000000001001000000; // D (0x0000000000000240) 
    12'h27e : LOC <=          63'b000000000000000000000000000000000000000000000000000001010000000; // D (0x0000000000000280) 
    12'hf43 : LOC <=          63'b000000000000000000000000000000000000000000000000000001100000000; // D (0x0000000000000300) 
    12'h695 : LOC <=          63'b000000000000000000000000000000000000000000000000000001000000000; // S (0x0000000000000200) 
//    12'hbbf : LOC <=          63'b000000000000000000000000000000000000000000000000000011000000000; // D (0x0000000000000600) 
//    12'h9f8 : LOC <=          63'b000000000000000000000000000000000000000000000000000101000000000; // D (0x0000000000000a00) 
//    12'hd76 : LOC <=          63'b000000000000000000000000000000000000000000000000001001000000000; // D (0x0000000000001200) 
//    12'h46a : LOC <=          63'b000000000000000000000000000000000000000000000000010001000000000; // D (0x0000000000002200) 
//    12'h36b : LOC <=          63'b000000000000000000000000000000000000000000000000100001000000000; // D (0x0000000000004200) 
//    12'hd69 : LOC <=          63'b000000000000000000000000000000000000000000000001000001000000000; // D (0x0000000000008200) 
//    12'h454 : LOC <=          63'b000000000000000000000000000000000000000000000010000001000000000; // D (0x0000000000010200) 
//    12'h317 : LOC <=          63'b000000000000000000000000000000000000000000000100000001000000000; // D (0x0000000000020200) 
//    12'hd91 : LOC <=          63'b000000000000000000000000000000000000000000001000000001000000000; // D (0x0000000000040200) 
//    12'h5a4 : LOC <=          63'b000000000000000000000000000000000000000000010000000001000000000; // D (0x0000000000080200) 
//    12'h0f7 : LOC <=          63'b000000000000000000000000000000000000000000100000000001000000000; // D (0x0000000000100200) 
//    12'ha51 : LOC <=          63'b000000000000000000000000000000000000000001000000000001000000000; // D (0x0000000000200200) 
//    12'ha24 : LOC <=          63'b000000000000000000000000000000000000000010000000000001000000000; // D (0x0000000000400200) 
//    12'hace : LOC <=          63'b000000000000000000000000000000000000000100000000000001000000000; // D (0x0000000000800200) 
//    12'hb1a : LOC <=          63'b000000000000000000000000000000000000001000000000000001000000000; // D (0x0000000001000200) 
//    12'h8b2 : LOC <=          63'b000000000000000000000000000000000000010000000000000001000000000; // D (0x0000000002000200) 
//    12'hfe2 : LOC <=          63'b000000000000000000000000000000000000100000000000000001000000000; // D (0x0000000004000200) 
//    12'h142 : LOC <=          63'b000000000000000000000000000000000001000000000000000001000000000; // D (0x0000000008000200) 
//    12'h93b : LOC <=          63'b000000000000000000000000000000000010000000000000000001000000000; // D (0x0000000010000200) 
//    12'hcf0 : LOC <=          63'b000000000000000000000000000000000100000000000000000001000000000; // D (0x0000000020000200) 
//    12'h766 : LOC <=          63'b000000000000000000000000000000001000000000000000000001000000000; // D (0x0000000040000200) 
//    12'h573 : LOC <=          63'b000000000000000000000000000000010000000000000000000001000000000; // D (0x0000000080000200) 
//    12'h159 : LOC <=          63'b000000000000000000000000000000100000000000000000000001000000000; // D (0x0000000100000200) 
//    12'h90d : LOC <=          63'b000000000000000000000000000001000000000000000000000001000000000; // D (0x0000000200000200) 
//    12'hc9c : LOC <=          63'b000000000000000000000000000010000000000000000000000001000000000; // D (0x0000000400000200) 
//    12'h7be : LOC <=          63'b000000000000000000000000000100000000000000000000000001000000000; // D (0x0000000800000200) 
//    12'h4c3 : LOC <=          63'b000000000000000000000000001000000000000000000000000001000000000; // D (0x0000001000000200) 
//    12'h239 : LOC <=          63'b000000000000000000000000010000000000000000000000000001000000000; // D (0x0000002000000200) 
//    12'hfcd : LOC <=          63'b000000000000000000000000100000000000000000000000000001000000000; // D (0x0000004000000200) 
//    12'h11c : LOC <=          63'b000000000000000000000001000000000000000000000000000001000000000; // D (0x0000008000000200) 
//    12'h987 : LOC <=          63'b000000000000000000000010000000000000000000000000000001000000000; // D (0x0000010000000200) 
//    12'hd88 : LOC <=          63'b000000000000000000000100000000000000000000000000000001000000000; // D (0x0000020000000200) 
//    12'h596 : LOC <=          63'b000000000000000000001000000000000000000000000000000001000000000; // D (0x0000040000000200) 
//    12'h093 : LOC <=          63'b000000000000000000010000000000000000000000000000000001000000000; // D (0x0000080000000200) 
//    12'ha99 : LOC <=          63'b000000000000000000100000000000000000000000000000000001000000000; // D (0x0000100000000200) 
//    12'hbb4 : LOC <=          63'b000000000000000001000000000000000000000000000000000001000000000; // D (0x0000200000000200) 
//    12'h9ee : LOC <=          63'b000000000000000010000000000000000000000000000000000001000000000; // D (0x0000400000000200) 
//    12'hd5a : LOC <=          63'b000000000000000100000000000000000000000000000000000001000000000; // D (0x0000800000000200) 
//    12'h432 : LOC <=          63'b000000000000001000000000000000000000000000000000000001000000000; // D (0x0001000000000200) 
//    12'h3db : LOC <=          63'b000000000000010000000000000000000000000000000000000001000000000; // D (0x0002000000000200) 
//    12'hc09 : LOC <=          63'b000000000000100000000000000000000000000000000000000001000000000; // D (0x0004000000000200) 
//    12'h694 : LOC <=          63'b000000000001000000000000000000000000000000000000000001000000000; // D (0x0008000000000200) 
//    12'h697 : LOC <=          63'b000000000010000000000000000000000000000000000000000001000000000; // D (0x0010000000000200) 
//    12'h691 : LOC <=          63'b000000000100000000000000000000000000000000000000000001000000000; // D (0x0020000000000200) 
//    12'h69d : LOC <=          63'b000000001000000000000000000000000000000000000000000001000000000; // D (0x0040000000000200) 
//    12'h685 : LOC <=          63'b000000010000000000000000000000000000000000000000000001000000000; // D (0x0080000000000200) 
//    12'h6b5 : LOC <=          63'b000000100000000000000000000000000000000000000000000001000000000; // D (0x0100000000000200) 
//    12'h6d5 : LOC <=          63'b000001000000000000000000000000000000000000000000000001000000000; // D (0x0200000000000200) 
//    12'h615 : LOC <=          63'b000010000000000000000000000000000000000000000000000001000000000; // D (0x0400000000000200) 
//    12'h795 : LOC <=          63'b000100000000000000000000000000000000000000000000000001000000000; // D (0x0800000000000200) 
//    12'h495 : LOC <=          63'b001000000000000000000000000000000000000000000000000001000000000; // D (0x1000000000000200) 
//    12'h295 : LOC <=          63'b010000000000000000000000000000000000000000000000000001000000000; // D (0x2000000000000200) 
//    12'he95 : LOC <=          63'b100000000000000000000000000000000000000000000000000001000000000; // D (0x4000000000000200) 
    12'h813 : LOC <=          63'b000000000000000000000000000000000000000000000000000010000000001; // D (0x0000000000000401) 
    12'h758 : LOC <=          63'b000000000000000000000000000000000000000000000000000010000000010; // D (0x0000000000000402) 
    12'hcf7 : LOC <=          63'b000000000000000000000000000000000000000000000000000010000000100; // D (0x0000000000000404) 
    12'he90 : LOC <=          63'b000000000000000000000000000000000000000000000000000010000001000; // D (0x0000000000000408) 
    12'ha5e : LOC <=          63'b000000000000000000000000000000000000000000000000000010000010000; // D (0x0000000000000410) 
    12'h3c2 : LOC <=          63'b000000000000000000000000000000000000000000000000000010000100000; // D (0x0000000000000420) 
    12'h5c3 : LOC <=          63'b000000000000000000000000000000000000000000000000000010001000000; // D (0x0000000000000440) 
    12'h9c1 : LOC <=          63'b000000000000000000000000000000000000000000000000000010010000000; // D (0x0000000000000480) 
    12'h4fc : LOC <=          63'b000000000000000000000000000000000000000000000000000010100000000; // D (0x0000000000000500) 
    12'hbbf : LOC <=          63'b000000000000000000000000000000000000000000000000000011000000000; // D (0x0000000000000600) 
    12'hd2a : LOC <=          63'b000000000000000000000000000000000000000000000000000010000000000; // S (0x0000000000000400) 
//    12'h247 : LOC <=          63'b000000000000000000000000000000000000000000000000000110000000000; // D (0x0000000000000c00) 
//    12'h6c9 : LOC <=          63'b000000000000000000000000000000000000000000000000001010000000000; // D (0x0000000000001400) 
//    12'hfd5 : LOC <=          63'b000000000000000000000000000000000000000000000000010010000000000; // D (0x0000000000002400) 
//    12'h8d4 : LOC <=          63'b000000000000000000000000000000000000000000000000100010000000000; // D (0x0000000000004400) 
//    12'h6d6 : LOC <=          63'b000000000000000000000000000000000000000000000001000010000000000; // D (0x0000000000008400) 
//    12'hfeb : LOC <=          63'b000000000000000000000000000000000000000000000010000010000000000; // D (0x0000000000010400) 
//    12'h8a8 : LOC <=          63'b000000000000000000000000000000000000000000000100000010000000000; // D (0x0000000000020400) 
//    12'h62e : LOC <=          63'b000000000000000000000000000000000000000000001000000010000000000; // D (0x0000000000040400) 
//    12'he1b : LOC <=          63'b000000000000000000000000000000000000000000010000000010000000000; // D (0x0000000000080400) 
//    12'hb48 : LOC <=          63'b000000000000000000000000000000000000000000100000000010000000000; // D (0x0000000000100400) 
//    12'h1ee : LOC <=          63'b000000000000000000000000000000000000000001000000000010000000000; // D (0x0000000000200400) 
//    12'h19b : LOC <=          63'b000000000000000000000000000000000000000010000000000010000000000; // D (0x0000000000400400) 
//    12'h171 : LOC <=          63'b000000000000000000000000000000000000000100000000000010000000000; // D (0x0000000000800400) 
//    12'h0a5 : LOC <=          63'b000000000000000000000000000000000000001000000000000010000000000; // D (0x0000000001000400) 
//    12'h30d : LOC <=          63'b000000000000000000000000000000000000010000000000000010000000000; // D (0x0000000002000400) 
//    12'h45d : LOC <=          63'b000000000000000000000000000000000000100000000000000010000000000; // D (0x0000000004000400) 
//    12'hafd : LOC <=          63'b000000000000000000000000000000000001000000000000000010000000000; // D (0x0000000008000400) 
//    12'h284 : LOC <=          63'b000000000000000000000000000000000010000000000000000010000000000; // D (0x0000000010000400) 
//    12'h74f : LOC <=          63'b000000000000000000000000000000000100000000000000000010000000000; // D (0x0000000020000400) 
//    12'hcd9 : LOC <=          63'b000000000000000000000000000000001000000000000000000010000000000; // D (0x0000000040000400) 
//    12'hecc : LOC <=          63'b000000000000000000000000000000010000000000000000000010000000000; // D (0x0000000080000400) 
//    12'hae6 : LOC <=          63'b000000000000000000000000000000100000000000000000000010000000000; // D (0x0000000100000400) 
//    12'h2b2 : LOC <=          63'b000000000000000000000000000001000000000000000000000010000000000; // D (0x0000000200000400) 
//    12'h723 : LOC <=          63'b000000000000000000000000000010000000000000000000000010000000000; // D (0x0000000400000400) 
//    12'hc01 : LOC <=          63'b000000000000000000000000000100000000000000000000000010000000000; // D (0x0000000800000400) 
//    12'hf7c : LOC <=          63'b000000000000000000000000001000000000000000000000000010000000000; // D (0x0000001000000400) 
//    12'h986 : LOC <=          63'b000000000000000000000000010000000000000000000000000010000000000; // D (0x0000002000000400) 
//    12'h472 : LOC <=          63'b000000000000000000000000100000000000000000000000000010000000000; // D (0x0000004000000400) 
//    12'haa3 : LOC <=          63'b000000000000000000000001000000000000000000000000000010000000000; // D (0x0000008000000400) 
//    12'h238 : LOC <=          63'b000000000000000000000010000000000000000000000000000010000000000; // D (0x0000010000000400) 
//    12'h637 : LOC <=          63'b000000000000000000000100000000000000000000000000000010000000000; // D (0x0000020000000400) 
//    12'he29 : LOC <=          63'b000000000000000000001000000000000000000000000000000010000000000; // D (0x0000040000000400) 
//    12'hb2c : LOC <=          63'b000000000000000000010000000000000000000000000000000010000000000; // D (0x0000080000000400) 
//    12'h126 : LOC <=          63'b000000000000000000100000000000000000000000000000000010000000000; // D (0x0000100000000400) 
//    12'h00b : LOC <=          63'b000000000000000001000000000000000000000000000000000010000000000; // D (0x0000200000000400) 
//    12'h251 : LOC <=          63'b000000000000000010000000000000000000000000000000000010000000000; // D (0x0000400000000400) 
//    12'h6e5 : LOC <=          63'b000000000000000100000000000000000000000000000000000010000000000; // D (0x0000800000000400) 
//    12'hf8d : LOC <=          63'b000000000000001000000000000000000000000000000000000010000000000; // D (0x0001000000000400) 
//    12'h864 : LOC <=          63'b000000000000010000000000000000000000000000000000000010000000000; // D (0x0002000000000400) 
//    12'h7b6 : LOC <=          63'b000000000000100000000000000000000000000000000000000010000000000; // D (0x0004000000000400) 
//    12'hd2b : LOC <=          63'b000000000001000000000000000000000000000000000000000010000000000; // D (0x0008000000000400) 
//    12'hd28 : LOC <=          63'b000000000010000000000000000000000000000000000000000010000000000; // D (0x0010000000000400) 
//    12'hd2e : LOC <=          63'b000000000100000000000000000000000000000000000000000010000000000; // D (0x0020000000000400) 
//    12'hd22 : LOC <=          63'b000000001000000000000000000000000000000000000000000010000000000; // D (0x0040000000000400) 
//    12'hd3a : LOC <=          63'b000000010000000000000000000000000000000000000000000010000000000; // D (0x0080000000000400) 
//    12'hd0a : LOC <=          63'b000000100000000000000000000000000000000000000000000010000000000; // D (0x0100000000000400) 
//    12'hd6a : LOC <=          63'b000001000000000000000000000000000000000000000000000010000000000; // D (0x0200000000000400) 
//    12'hdaa : LOC <=          63'b000010000000000000000000000000000000000000000000000010000000000; // D (0x0400000000000400) 
//    12'hc2a : LOC <=          63'b000100000000000000000000000000000000000000000000000010000000000; // D (0x0800000000000400) 
//    12'hf2a : LOC <=          63'b001000000000000000000000000000000000000000000000000010000000000; // D (0x1000000000000400) 
//    12'h92a : LOC <=          63'b010000000000000000000000000000000000000000000000000010000000000; // D (0x2000000000000400) 
//    12'h52a : LOC <=          63'b100000000000000000000000000000000000000000000000000010000000000; // D (0x4000000000000400) 
    12'ha54 : LOC <=          63'b000000000000000000000000000000000000000000000000000100000000001; // D (0x0000000000000801) 
    12'h51f : LOC <=          63'b000000000000000000000000000000000000000000000000000100000000010; // D (0x0000000000000802) 
    12'heb0 : LOC <=          63'b000000000000000000000000000000000000000000000000000100000000100; // D (0x0000000000000804) 
    12'hcd7 : LOC <=          63'b000000000000000000000000000000000000000000000000000100000001000; // D (0x0000000000000808) 
    12'h819 : LOC <=          63'b000000000000000000000000000000000000000000000000000100000010000; // D (0x0000000000000810) 
    12'h185 : LOC <=          63'b000000000000000000000000000000000000000000000000000100000100000; // D (0x0000000000000820) 
    12'h784 : LOC <=          63'b000000000000000000000000000000000000000000000000000100001000000; // D (0x0000000000000840) 
    12'hb86 : LOC <=          63'b000000000000000000000000000000000000000000000000000100010000000; // D (0x0000000000000880) 
    12'h6bb : LOC <=          63'b000000000000000000000000000000000000000000000000000100100000000; // D (0x0000000000000900) 
    12'h9f8 : LOC <=          63'b000000000000000000000000000000000000000000000000000101000000000; // D (0x0000000000000a00) 
    12'h247 : LOC <=          63'b000000000000000000000000000000000000000000000000000110000000000; // D (0x0000000000000c00) 
    12'hf6d : LOC <=          63'b000000000000000000000000000000000000000000000000000100000000000; // S (0x0000000000000800) 
//    12'h48e : LOC <=          63'b000000000000000000000000000000000000000000000000001100000000000; // D (0x0000000000001800) 
//    12'hd92 : LOC <=          63'b000000000000000000000000000000000000000000000000010100000000000; // D (0x0000000000002800) 
//    12'ha93 : LOC <=          63'b000000000000000000000000000000000000000000000000100100000000000; // D (0x0000000000004800) 
//    12'h491 : LOC <=          63'b000000000000000000000000000000000000000000000001000100000000000; // D (0x0000000000008800) 
//    12'hdac : LOC <=          63'b000000000000000000000000000000000000000000000010000100000000000; // D (0x0000000000010800) 
//    12'haef : LOC <=          63'b000000000000000000000000000000000000000000000100000100000000000; // D (0x0000000000020800) 
//    12'h469 : LOC <=          63'b000000000000000000000000000000000000000000001000000100000000000; // D (0x0000000000040800) 
//    12'hc5c : LOC <=          63'b000000000000000000000000000000000000000000010000000100000000000; // D (0x0000000000080800) 
//    12'h90f : LOC <=          63'b000000000000000000000000000000000000000000100000000100000000000; // D (0x0000000000100800) 
//    12'h3a9 : LOC <=          63'b000000000000000000000000000000000000000001000000000100000000000; // D (0x0000000000200800) 
//    12'h3dc : LOC <=          63'b000000000000000000000000000000000000000010000000000100000000000; // D (0x0000000000400800) 
//    12'h336 : LOC <=          63'b000000000000000000000000000000000000000100000000000100000000000; // D (0x0000000000800800) 
//    12'h2e2 : LOC <=          63'b000000000000000000000000000000000000001000000000000100000000000; // D (0x0000000001000800) 
//    12'h14a : LOC <=          63'b000000000000000000000000000000000000010000000000000100000000000; // D (0x0000000002000800) 
//    12'h61a : LOC <=          63'b000000000000000000000000000000000000100000000000000100000000000; // D (0x0000000004000800) 
//    12'h8ba : LOC <=          63'b000000000000000000000000000000000001000000000000000100000000000; // D (0x0000000008000800) 
//    12'h0c3 : LOC <=          63'b000000000000000000000000000000000010000000000000000100000000000; // D (0x0000000010000800) 
//    12'h508 : LOC <=          63'b000000000000000000000000000000000100000000000000000100000000000; // D (0x0000000020000800) 
//    12'he9e : LOC <=          63'b000000000000000000000000000000001000000000000000000100000000000; // D (0x0000000040000800) 
//    12'hc8b : LOC <=          63'b000000000000000000000000000000010000000000000000000100000000000; // D (0x0000000080000800) 
//    12'h8a1 : LOC <=          63'b000000000000000000000000000000100000000000000000000100000000000; // D (0x0000000100000800) 
//    12'h0f5 : LOC <=          63'b000000000000000000000000000001000000000000000000000100000000000; // D (0x0000000200000800) 
//    12'h564 : LOC <=          63'b000000000000000000000000000010000000000000000000000100000000000; // D (0x0000000400000800) 
//    12'he46 : LOC <=          63'b000000000000000000000000000100000000000000000000000100000000000; // D (0x0000000800000800) 
//    12'hd3b : LOC <=          63'b000000000000000000000000001000000000000000000000000100000000000; // D (0x0000001000000800) 
//    12'hbc1 : LOC <=          63'b000000000000000000000000010000000000000000000000000100000000000; // D (0x0000002000000800) 
//    12'h635 : LOC <=          63'b000000000000000000000000100000000000000000000000000100000000000; // D (0x0000004000000800) 
//    12'h8e4 : LOC <=          63'b000000000000000000000001000000000000000000000000000100000000000; // D (0x0000008000000800) 
//    12'h07f : LOC <=          63'b000000000000000000000010000000000000000000000000000100000000000; // D (0x0000010000000800) 
//    12'h470 : LOC <=          63'b000000000000000000000100000000000000000000000000000100000000000; // D (0x0000020000000800) 
//    12'hc6e : LOC <=          63'b000000000000000000001000000000000000000000000000000100000000000; // D (0x0000040000000800) 
//    12'h96b : LOC <=          63'b000000000000000000010000000000000000000000000000000100000000000; // D (0x0000080000000800) 
//    12'h361 : LOC <=          63'b000000000000000000100000000000000000000000000000000100000000000; // D (0x0000100000000800) 
//    12'h24c : LOC <=          63'b000000000000000001000000000000000000000000000000000100000000000; // D (0x0000200000000800) 
//    12'h016 : LOC <=          63'b000000000000000010000000000000000000000000000000000100000000000; // D (0x0000400000000800) 
//    12'h4a2 : LOC <=          63'b000000000000000100000000000000000000000000000000000100000000000; // D (0x0000800000000800) 
//    12'hdca : LOC <=          63'b000000000000001000000000000000000000000000000000000100000000000; // D (0x0001000000000800) 
//    12'ha23 : LOC <=          63'b000000000000010000000000000000000000000000000000000100000000000; // D (0x0002000000000800) 
//    12'h5f1 : LOC <=          63'b000000000000100000000000000000000000000000000000000100000000000; // D (0x0004000000000800) 
//    12'hf6c : LOC <=          63'b000000000001000000000000000000000000000000000000000100000000000; // D (0x0008000000000800) 
//    12'hf6f : LOC <=          63'b000000000010000000000000000000000000000000000000000100000000000; // D (0x0010000000000800) 
//    12'hf69 : LOC <=          63'b000000000100000000000000000000000000000000000000000100000000000; // D (0x0020000000000800) 
//    12'hf65 : LOC <=          63'b000000001000000000000000000000000000000000000000000100000000000; // D (0x0040000000000800) 
//    12'hf7d : LOC <=          63'b000000010000000000000000000000000000000000000000000100000000000; // D (0x0080000000000800) 
//    12'hf4d : LOC <=          63'b000000100000000000000000000000000000000000000000000100000000000; // D (0x0100000000000800) 
//    12'hf2d : LOC <=          63'b000001000000000000000000000000000000000000000000000100000000000; // D (0x0200000000000800) 
//    12'hfed : LOC <=          63'b000010000000000000000000000000000000000000000000000100000000000; // D (0x0400000000000800) 
//    12'he6d : LOC <=          63'b000100000000000000000000000000000000000000000000000100000000000; // D (0x0800000000000800) 
//    12'hd6d : LOC <=          63'b001000000000000000000000000000000000000000000000000100000000000; // D (0x1000000000000800) 
//    12'hb6d : LOC <=          63'b010000000000000000000000000000000000000000000000000100000000000; // D (0x2000000000000800) 
//    12'h76d : LOC <=          63'b100000000000000000000000000000000000000000000000000100000000000; // D (0x4000000000000800) 
    12'heda : LOC <=          63'b000000000000000000000000000000000000000000000000001000000000001; // D (0x0000000000001001) 
    12'h191 : LOC <=          63'b000000000000000000000000000000000000000000000000001000000000010; // D (0x0000000000001002) 
    12'ha3e : LOC <=          63'b000000000000000000000000000000000000000000000000001000000000100; // D (0x0000000000001004) 
    12'h859 : LOC <=          63'b000000000000000000000000000000000000000000000000001000000001000; // D (0x0000000000001008) 
    12'hc97 : LOC <=          63'b000000000000000000000000000000000000000000000000001000000010000; // D (0x0000000000001010) 
    12'h50b : LOC <=          63'b000000000000000000000000000000000000000000000000001000000100000; // D (0x0000000000001020) 
    12'h30a : LOC <=          63'b000000000000000000000000000000000000000000000000001000001000000; // D (0x0000000000001040) 
    12'hf08 : LOC <=          63'b000000000000000000000000000000000000000000000000001000010000000; // D (0x0000000000001080) 
    12'h235 : LOC <=          63'b000000000000000000000000000000000000000000000000001000100000000; // D (0x0000000000001100) 
    12'hd76 : LOC <=          63'b000000000000000000000000000000000000000000000000001001000000000; // D (0x0000000000001200) 
    12'h6c9 : LOC <=          63'b000000000000000000000000000000000000000000000000001010000000000; // D (0x0000000000001400) 
    12'h48e : LOC <=          63'b000000000000000000000000000000000000000000000000001100000000000; // D (0x0000000000001800) 
    12'hbe3 : LOC <=          63'b000000000000000000000000000000000000000000000000001000000000000; // S (0x0000000000001000) 
//    12'h91c : LOC <=          63'b000000000000000000000000000000000000000000000000011000000000000; // D (0x0000000000003000) 
//    12'he1d : LOC <=          63'b000000000000000000000000000000000000000000000000101000000000000; // D (0x0000000000005000) 
//    12'h01f : LOC <=          63'b000000000000000000000000000000000000000000000001001000000000000; // D (0x0000000000009000) 
//    12'h922 : LOC <=          63'b000000000000000000000000000000000000000000000010001000000000000; // D (0x0000000000011000) 
//    12'he61 : LOC <=          63'b000000000000000000000000000000000000000000000100001000000000000; // D (0x0000000000021000) 
//    12'h0e7 : LOC <=          63'b000000000000000000000000000000000000000000001000001000000000000; // D (0x0000000000041000) 
//    12'h8d2 : LOC <=          63'b000000000000000000000000000000000000000000010000001000000000000; // D (0x0000000000081000) 
//    12'hd81 : LOC <=          63'b000000000000000000000000000000000000000000100000001000000000000; // D (0x0000000000101000) 
//    12'h727 : LOC <=          63'b000000000000000000000000000000000000000001000000001000000000000; // D (0x0000000000201000) 
//    12'h752 : LOC <=          63'b000000000000000000000000000000000000000010000000001000000000000; // D (0x0000000000401000) 
//    12'h7b8 : LOC <=          63'b000000000000000000000000000000000000000100000000001000000000000; // D (0x0000000000801000) 
//    12'h66c : LOC <=          63'b000000000000000000000000000000000000001000000000001000000000000; // D (0x0000000001001000) 
//    12'h5c4 : LOC <=          63'b000000000000000000000000000000000000010000000000001000000000000; // D (0x0000000002001000) 
//    12'h294 : LOC <=          63'b000000000000000000000000000000000000100000000000001000000000000; // D (0x0000000004001000) 
//    12'hc34 : LOC <=          63'b000000000000000000000000000000000001000000000000001000000000000; // D (0x0000000008001000) 
//    12'h44d : LOC <=          63'b000000000000000000000000000000000010000000000000001000000000000; // D (0x0000000010001000) 
//    12'h186 : LOC <=          63'b000000000000000000000000000000000100000000000000001000000000000; // D (0x0000000020001000) 
//    12'ha10 : LOC <=          63'b000000000000000000000000000000001000000000000000001000000000000; // D (0x0000000040001000) 
//    12'h805 : LOC <=          63'b000000000000000000000000000000010000000000000000001000000000000; // D (0x0000000080001000) 
//    12'hc2f : LOC <=          63'b000000000000000000000000000000100000000000000000001000000000000; // D (0x0000000100001000) 
//    12'h47b : LOC <=          63'b000000000000000000000000000001000000000000000000001000000000000; // D (0x0000000200001000) 
//    12'h1ea : LOC <=          63'b000000000000000000000000000010000000000000000000001000000000000; // D (0x0000000400001000) 
//    12'hac8 : LOC <=          63'b000000000000000000000000000100000000000000000000001000000000000; // D (0x0000000800001000) 
//    12'h9b5 : LOC <=          63'b000000000000000000000000001000000000000000000000001000000000000; // D (0x0000001000001000) 
//    12'hf4f : LOC <=          63'b000000000000000000000000010000000000000000000000001000000000000; // D (0x0000002000001000) 
//    12'h2bb : LOC <=          63'b000000000000000000000000100000000000000000000000001000000000000; // D (0x0000004000001000) 
//    12'hc6a : LOC <=          63'b000000000000000000000001000000000000000000000000001000000000000; // D (0x0000008000001000) 
//    12'h4f1 : LOC <=          63'b000000000000000000000010000000000000000000000000001000000000000; // D (0x0000010000001000) 
//    12'h0fe : LOC <=          63'b000000000000000000000100000000000000000000000000001000000000000; // D (0x0000020000001000) 
//    12'h8e0 : LOC <=          63'b000000000000000000001000000000000000000000000000001000000000000; // D (0x0000040000001000) 
//    12'hde5 : LOC <=          63'b000000000000000000010000000000000000000000000000001000000000000; // D (0x0000080000001000) 
//    12'h7ef : LOC <=          63'b000000000000000000100000000000000000000000000000001000000000000; // D (0x0000100000001000) 
//    12'h6c2 : LOC <=          63'b000000000000000001000000000000000000000000000000001000000000000; // D (0x0000200000001000) 
//    12'h498 : LOC <=          63'b000000000000000010000000000000000000000000000000001000000000000; // D (0x0000400000001000) 
//    12'h02c : LOC <=          63'b000000000000000100000000000000000000000000000000001000000000000; // D (0x0000800000001000) 
//    12'h944 : LOC <=          63'b000000000000001000000000000000000000000000000000001000000000000; // D (0x0001000000001000) 
//    12'head : LOC <=          63'b000000000000010000000000000000000000000000000000001000000000000; // D (0x0002000000001000) 
//    12'h17f : LOC <=          63'b000000000000100000000000000000000000000000000000001000000000000; // D (0x0004000000001000) 
//    12'hbe2 : LOC <=          63'b000000000001000000000000000000000000000000000000001000000000000; // D (0x0008000000001000) 
//    12'hbe1 : LOC <=          63'b000000000010000000000000000000000000000000000000001000000000000; // D (0x0010000000001000) 
//    12'hbe7 : LOC <=          63'b000000000100000000000000000000000000000000000000001000000000000; // D (0x0020000000001000) 
//    12'hbeb : LOC <=          63'b000000001000000000000000000000000000000000000000001000000000000; // D (0x0040000000001000) 
//    12'hbf3 : LOC <=          63'b000000010000000000000000000000000000000000000000001000000000000; // D (0x0080000000001000) 
//    12'hbc3 : LOC <=          63'b000000100000000000000000000000000000000000000000001000000000000; // D (0x0100000000001000) 
//    12'hba3 : LOC <=          63'b000001000000000000000000000000000000000000000000001000000000000; // D (0x0200000000001000) 
//    12'hb63 : LOC <=          63'b000010000000000000000000000000000000000000000000001000000000000; // D (0x0400000000001000) 
//    12'hae3 : LOC <=          63'b000100000000000000000000000000000000000000000000001000000000000; // D (0x0800000000001000) 
//    12'h9e3 : LOC <=          63'b001000000000000000000000000000000000000000000000001000000000000; // D (0x1000000000001000) 
//    12'hfe3 : LOC <=          63'b010000000000000000000000000000000000000000000000001000000000000; // D (0x2000000000001000) 
//    12'h3e3 : LOC <=          63'b100000000000000000000000000000000000000000000000001000000000000; // D (0x4000000000001000) 
    12'h7c6 : LOC <=          63'b000000000000000000000000000000000000000000000000010000000000001; // D (0x0000000000002001) 
    12'h88d : LOC <=          63'b000000000000000000000000000000000000000000000000010000000000010; // D (0x0000000000002002) 
    12'h322 : LOC <=          63'b000000000000000000000000000000000000000000000000010000000000100; // D (0x0000000000002004) 
    12'h145 : LOC <=          63'b000000000000000000000000000000000000000000000000010000000001000; // D (0x0000000000002008) 
    12'h58b : LOC <=          63'b000000000000000000000000000000000000000000000000010000000010000; // D (0x0000000000002010) 
    12'hc17 : LOC <=          63'b000000000000000000000000000000000000000000000000010000000100000; // D (0x0000000000002020) 
    12'ha16 : LOC <=          63'b000000000000000000000000000000000000000000000000010000001000000; // D (0x0000000000002040) 
    12'h614 : LOC <=          63'b000000000000000000000000000000000000000000000000010000010000000; // D (0x0000000000002080) 
    12'hb29 : LOC <=          63'b000000000000000000000000000000000000000000000000010000100000000; // D (0x0000000000002100) 
    12'h46a : LOC <=          63'b000000000000000000000000000000000000000000000000010001000000000; // D (0x0000000000002200) 
    12'hfd5 : LOC <=          63'b000000000000000000000000000000000000000000000000010010000000000; // D (0x0000000000002400) 
    12'hd92 : LOC <=          63'b000000000000000000000000000000000000000000000000010100000000000; // D (0x0000000000002800) 
    12'h91c : LOC <=          63'b000000000000000000000000000000000000000000000000011000000000000; // D (0x0000000000003000) 
    12'h2ff : LOC <=          63'b000000000000000000000000000000000000000000000000010000000000000; // S (0x0000000000002000) 
//    12'h701 : LOC <=          63'b000000000000000000000000000000000000000000000000110000000000000; // D (0x0000000000006000) 
//    12'h903 : LOC <=          63'b000000000000000000000000000000000000000000000001010000000000000; // D (0x000000000000a000) 
//    12'h03e : LOC <=          63'b000000000000000000000000000000000000000000000010010000000000000; // D (0x0000000000012000) 
//    12'h77d : LOC <=          63'b000000000000000000000000000000000000000000000100010000000000000; // D (0x0000000000022000) 
//    12'h9fb : LOC <=          63'b000000000000000000000000000000000000000000001000010000000000000; // D (0x0000000000042000) 
//    12'h1ce : LOC <=          63'b000000000000000000000000000000000000000000010000010000000000000; // D (0x0000000000082000) 
//    12'h49d : LOC <=          63'b000000000000000000000000000000000000000000100000010000000000000; // D (0x0000000000102000) 
//    12'he3b : LOC <=          63'b000000000000000000000000000000000000000001000000010000000000000; // D (0x0000000000202000) 
//    12'he4e : LOC <=          63'b000000000000000000000000000000000000000010000000010000000000000; // D (0x0000000000402000) 
//    12'hea4 : LOC <=          63'b000000000000000000000000000000000000000100000000010000000000000; // D (0x0000000000802000) 
//    12'hf70 : LOC <=          63'b000000000000000000000000000000000000001000000000010000000000000; // D (0x0000000001002000) 
//    12'hcd8 : LOC <=          63'b000000000000000000000000000000000000010000000000010000000000000; // D (0x0000000002002000) 
//    12'hb88 : LOC <=          63'b000000000000000000000000000000000000100000000000010000000000000; // D (0x0000000004002000) 
//    12'h528 : LOC <=          63'b000000000000000000000000000000000001000000000000010000000000000; // D (0x0000000008002000) 
//    12'hd51 : LOC <=          63'b000000000000000000000000000000000010000000000000010000000000000; // D (0x0000000010002000) 
//    12'h89a : LOC <=          63'b000000000000000000000000000000000100000000000000010000000000000; // D (0x0000000020002000) 
//    12'h30c : LOC <=          63'b000000000000000000000000000000001000000000000000010000000000000; // D (0x0000000040002000) 
//    12'h119 : LOC <=          63'b000000000000000000000000000000010000000000000000010000000000000; // D (0x0000000080002000) 
//    12'h533 : LOC <=          63'b000000000000000000000000000000100000000000000000010000000000000; // D (0x0000000100002000) 
//    12'hd67 : LOC <=          63'b000000000000000000000000000001000000000000000000010000000000000; // D (0x0000000200002000) 
//    12'h8f6 : LOC <=          63'b000000000000000000000000000010000000000000000000010000000000000; // D (0x0000000400002000) 
//    12'h3d4 : LOC <=          63'b000000000000000000000000000100000000000000000000010000000000000; // D (0x0000000800002000) 
//    12'h0a9 : LOC <=          63'b000000000000000000000000001000000000000000000000010000000000000; // D (0x0000001000002000) 
//    12'h653 : LOC <=          63'b000000000000000000000000010000000000000000000000010000000000000; // D (0x0000002000002000) 
//    12'hba7 : LOC <=          63'b000000000000000000000000100000000000000000000000010000000000000; // D (0x0000004000002000) 
//    12'h576 : LOC <=          63'b000000000000000000000001000000000000000000000000010000000000000; // D (0x0000008000002000) 
//    12'hded : LOC <=          63'b000000000000000000000010000000000000000000000000010000000000000; // D (0x0000010000002000) 
//    12'h9e2 : LOC <=          63'b000000000000000000000100000000000000000000000000010000000000000; // D (0x0000020000002000) 
//    12'h1fc : LOC <=          63'b000000000000000000001000000000000000000000000000010000000000000; // D (0x0000040000002000) 
//    12'h4f9 : LOC <=          63'b000000000000000000010000000000000000000000000000010000000000000; // D (0x0000080000002000) 
//    12'hef3 : LOC <=          63'b000000000000000000100000000000000000000000000000010000000000000; // D (0x0000100000002000) 
//    12'hfde : LOC <=          63'b000000000000000001000000000000000000000000000000010000000000000; // D (0x0000200000002000) 
//    12'hd84 : LOC <=          63'b000000000000000010000000000000000000000000000000010000000000000; // D (0x0000400000002000) 
//    12'h930 : LOC <=          63'b000000000000000100000000000000000000000000000000010000000000000; // D (0x0000800000002000) 
//    12'h058 : LOC <=          63'b000000000000001000000000000000000000000000000000010000000000000; // D (0x0001000000002000) 
//    12'h7b1 : LOC <=          63'b000000000000010000000000000000000000000000000000010000000000000; // D (0x0002000000002000) 
//    12'h863 : LOC <=          63'b000000000000100000000000000000000000000000000000010000000000000; // D (0x0004000000002000) 
//    12'h2fe : LOC <=          63'b000000000001000000000000000000000000000000000000010000000000000; // D (0x0008000000002000) 
//    12'h2fd : LOC <=          63'b000000000010000000000000000000000000000000000000010000000000000; // D (0x0010000000002000) 
//    12'h2fb : LOC <=          63'b000000000100000000000000000000000000000000000000010000000000000; // D (0x0020000000002000) 
//    12'h2f7 : LOC <=          63'b000000001000000000000000000000000000000000000000010000000000000; // D (0x0040000000002000) 
//    12'h2ef : LOC <=          63'b000000010000000000000000000000000000000000000000010000000000000; // D (0x0080000000002000) 
//    12'h2df : LOC <=          63'b000000100000000000000000000000000000000000000000010000000000000; // D (0x0100000000002000) 
//    12'h2bf : LOC <=          63'b000001000000000000000000000000000000000000000000010000000000000; // D (0x0200000000002000) 
//    12'h27f : LOC <=          63'b000010000000000000000000000000000000000000000000010000000000000; // D (0x0400000000002000) 
//    12'h3ff : LOC <=          63'b000100000000000000000000000000000000000000000000010000000000000; // D (0x0800000000002000) 
//    12'h0ff : LOC <=          63'b001000000000000000000000000000000000000000000000010000000000000; // D (0x1000000000002000) 
//    12'h6ff : LOC <=          63'b010000000000000000000000000000000000000000000000010000000000000; // D (0x2000000000002000) 
//    12'haff : LOC <=          63'b100000000000000000000000000000000000000000000000010000000000000; // D (0x4000000000002000) 
    12'h0c7 : LOC <=          63'b000000000000000000000000000000000000000000000000100000000000001; // D (0x0000000000004001) 
    12'hf8c : LOC <=          63'b000000000000000000000000000000000000000000000000100000000000010; // D (0x0000000000004002) 
    12'h423 : LOC <=          63'b000000000000000000000000000000000000000000000000100000000000100; // D (0x0000000000004004) 
    12'h644 : LOC <=          63'b000000000000000000000000000000000000000000000000100000000001000; // D (0x0000000000004008) 
    12'h28a : LOC <=          63'b000000000000000000000000000000000000000000000000100000000010000; // D (0x0000000000004010) 
    12'hb16 : LOC <=          63'b000000000000000000000000000000000000000000000000100000000100000; // D (0x0000000000004020) 
    12'hd17 : LOC <=          63'b000000000000000000000000000000000000000000000000100000001000000; // D (0x0000000000004040) 
    12'h115 : LOC <=          63'b000000000000000000000000000000000000000000000000100000010000000; // D (0x0000000000004080) 
    12'hc28 : LOC <=          63'b000000000000000000000000000000000000000000000000100000100000000; // D (0x0000000000004100) 
    12'h36b : LOC <=          63'b000000000000000000000000000000000000000000000000100001000000000; // D (0x0000000000004200) 
    12'h8d4 : LOC <=          63'b000000000000000000000000000000000000000000000000100010000000000; // D (0x0000000000004400) 
    12'ha93 : LOC <=          63'b000000000000000000000000000000000000000000000000100100000000000; // D (0x0000000000004800) 
    12'he1d : LOC <=          63'b000000000000000000000000000000000000000000000000101000000000000; // D (0x0000000000005000) 
    12'h701 : LOC <=          63'b000000000000000000000000000000000000000000000000110000000000000; // D (0x0000000000006000) 
    12'h5fe : LOC <=          63'b000000000000000000000000000000000000000000000000100000000000000; // S (0x0000000000004000) 
//    12'he02 : LOC <=          63'b000000000000000000000000000000000000000000000001100000000000000; // D (0x000000000000c000) 
//    12'h73f : LOC <=          63'b000000000000000000000000000000000000000000000010100000000000000; // D (0x0000000000014000) 
//    12'h07c : LOC <=          63'b000000000000000000000000000000000000000000000100100000000000000; // D (0x0000000000024000) 
//    12'hefa : LOC <=          63'b000000000000000000000000000000000000000000001000100000000000000; // D (0x0000000000044000) 
//    12'h6cf : LOC <=          63'b000000000000000000000000000000000000000000010000100000000000000; // D (0x0000000000084000) 
//    12'h39c : LOC <=          63'b000000000000000000000000000000000000000000100000100000000000000; // D (0x0000000000104000) 
//    12'h93a : LOC <=          63'b000000000000000000000000000000000000000001000000100000000000000; // D (0x0000000000204000) 
//    12'h94f : LOC <=          63'b000000000000000000000000000000000000000010000000100000000000000; // D (0x0000000000404000) 
//    12'h9a5 : LOC <=          63'b000000000000000000000000000000000000000100000000100000000000000; // D (0x0000000000804000) 
//    12'h871 : LOC <=          63'b000000000000000000000000000000000000001000000000100000000000000; // D (0x0000000001004000) 
//    12'hbd9 : LOC <=          63'b000000000000000000000000000000000000010000000000100000000000000; // D (0x0000000002004000) 
//    12'hc89 : LOC <=          63'b000000000000000000000000000000000000100000000000100000000000000; // D (0x0000000004004000) 
//    12'h229 : LOC <=          63'b000000000000000000000000000000000001000000000000100000000000000; // D (0x0000000008004000) 
//    12'ha50 : LOC <=          63'b000000000000000000000000000000000010000000000000100000000000000; // D (0x0000000010004000) 
//    12'hf9b : LOC <=          63'b000000000000000000000000000000000100000000000000100000000000000; // D (0x0000000020004000) 
//    12'h40d : LOC <=          63'b000000000000000000000000000000001000000000000000100000000000000; // D (0x0000000040004000) 
//    12'h618 : LOC <=          63'b000000000000000000000000000000010000000000000000100000000000000; // D (0x0000000080004000) 
//    12'h232 : LOC <=          63'b000000000000000000000000000000100000000000000000100000000000000; // D (0x0000000100004000) 
//    12'ha66 : LOC <=          63'b000000000000000000000000000001000000000000000000100000000000000; // D (0x0000000200004000) 
//    12'hff7 : LOC <=          63'b000000000000000000000000000010000000000000000000100000000000000; // D (0x0000000400004000) 
//    12'h4d5 : LOC <=          63'b000000000000000000000000000100000000000000000000100000000000000; // D (0x0000000800004000) 
//    12'h7a8 : LOC <=          63'b000000000000000000000000001000000000000000000000100000000000000; // D (0x0000001000004000) 
//    12'h152 : LOC <=          63'b000000000000000000000000010000000000000000000000100000000000000; // D (0x0000002000004000) 
//    12'hca6 : LOC <=          63'b000000000000000000000000100000000000000000000000100000000000000; // D (0x0000004000004000) 
//    12'h277 : LOC <=          63'b000000000000000000000001000000000000000000000000100000000000000; // D (0x0000008000004000) 
//    12'haec : LOC <=          63'b000000000000000000000010000000000000000000000000100000000000000; // D (0x0000010000004000) 
//    12'hee3 : LOC <=          63'b000000000000000000000100000000000000000000000000100000000000000; // D (0x0000020000004000) 
//    12'h6fd : LOC <=          63'b000000000000000000001000000000000000000000000000100000000000000; // D (0x0000040000004000) 
//    12'h3f8 : LOC <=          63'b000000000000000000010000000000000000000000000000100000000000000; // D (0x0000080000004000) 
//    12'h9f2 : LOC <=          63'b000000000000000000100000000000000000000000000000100000000000000; // D (0x0000100000004000) 
//    12'h8df : LOC <=          63'b000000000000000001000000000000000000000000000000100000000000000; // D (0x0000200000004000) 
//    12'ha85 : LOC <=          63'b000000000000000010000000000000000000000000000000100000000000000; // D (0x0000400000004000) 
//    12'he31 : LOC <=          63'b000000000000000100000000000000000000000000000000100000000000000; // D (0x0000800000004000) 
//    12'h759 : LOC <=          63'b000000000000001000000000000000000000000000000000100000000000000; // D (0x0001000000004000) 
//    12'h0b0 : LOC <=          63'b000000000000010000000000000000000000000000000000100000000000000; // D (0x0002000000004000) 
//    12'hf62 : LOC <=          63'b000000000000100000000000000000000000000000000000100000000000000; // D (0x0004000000004000) 
//    12'h5ff : LOC <=          63'b000000000001000000000000000000000000000000000000100000000000000; // D (0x0008000000004000) 
//    12'h5fc : LOC <=          63'b000000000010000000000000000000000000000000000000100000000000000; // D (0x0010000000004000) 
//    12'h5fa : LOC <=          63'b000000000100000000000000000000000000000000000000100000000000000; // D (0x0020000000004000) 
//    12'h5f6 : LOC <=          63'b000000001000000000000000000000000000000000000000100000000000000; // D (0x0040000000004000) 
//    12'h5ee : LOC <=          63'b000000010000000000000000000000000000000000000000100000000000000; // D (0x0080000000004000) 
//    12'h5de : LOC <=          63'b000000100000000000000000000000000000000000000000100000000000000; // D (0x0100000000004000) 
//    12'h5be : LOC <=          63'b000001000000000000000000000000000000000000000000100000000000000; // D (0x0200000000004000) 
//    12'h57e : LOC <=          63'b000010000000000000000000000000000000000000000000100000000000000; // D (0x0400000000004000) 
//    12'h4fe : LOC <=          63'b000100000000000000000000000000000000000000000000100000000000000; // D (0x0800000000004000) 
//    12'h7fe : LOC <=          63'b001000000000000000000000000000000000000000000000100000000000000; // D (0x1000000000004000) 
//    12'h1fe : LOC <=          63'b010000000000000000000000000000000000000000000000100000000000000; // D (0x2000000000004000) 
//    12'hdfe : LOC <=          63'b100000000000000000000000000000000000000000000000100000000000000; // D (0x4000000000004000) 
    12'hec5 : LOC <=          63'b000000000000000000000000000000000000000000000001000000000000001; // D (0x0000000000008001) 
    12'h18e : LOC <=          63'b000000000000000000000000000000000000000000000001000000000000010; // D (0x0000000000008002) 
    12'ha21 : LOC <=          63'b000000000000000000000000000000000000000000000001000000000000100; // D (0x0000000000008004) 
    12'h846 : LOC <=          63'b000000000000000000000000000000000000000000000001000000000001000; // D (0x0000000000008008) 
    12'hc88 : LOC <=          63'b000000000000000000000000000000000000000000000001000000000010000; // D (0x0000000000008010) 
    12'h514 : LOC <=          63'b000000000000000000000000000000000000000000000001000000000100000; // D (0x0000000000008020) 
    12'h315 : LOC <=          63'b000000000000000000000000000000000000000000000001000000001000000; // D (0x0000000000008040) 
    12'hf17 : LOC <=          63'b000000000000000000000000000000000000000000000001000000010000000; // D (0x0000000000008080) 
    12'h22a : LOC <=          63'b000000000000000000000000000000000000000000000001000000100000000; // D (0x0000000000008100) 
    12'hd69 : LOC <=          63'b000000000000000000000000000000000000000000000001000001000000000; // D (0x0000000000008200) 
    12'h6d6 : LOC <=          63'b000000000000000000000000000000000000000000000001000010000000000; // D (0x0000000000008400) 
    12'h491 : LOC <=          63'b000000000000000000000000000000000000000000000001000100000000000; // D (0x0000000000008800) 
    12'h01f : LOC <=          63'b000000000000000000000000000000000000000000000001001000000000000; // D (0x0000000000009000) 
    12'h903 : LOC <=          63'b000000000000000000000000000000000000000000000001010000000000000; // D (0x000000000000a000) 
    12'he02 : LOC <=          63'b000000000000000000000000000000000000000000000001100000000000000; // D (0x000000000000c000) 
    12'hbfc : LOC <=          63'b000000000000000000000000000000000000000000000001000000000000000; // S (0x0000000000008000) 
//    12'h93d : LOC <=          63'b000000000000000000000000000000000000000000000011000000000000000; // D (0x0000000000018000) 
//    12'he7e : LOC <=          63'b000000000000000000000000000000000000000000000101000000000000000; // D (0x0000000000028000) 
//    12'h0f8 : LOC <=          63'b000000000000000000000000000000000000000000001001000000000000000; // D (0x0000000000048000) 
//    12'h8cd : LOC <=          63'b000000000000000000000000000000000000000000010001000000000000000; // D (0x0000000000088000) 
//    12'hd9e : LOC <=          63'b000000000000000000000000000000000000000000100001000000000000000; // D (0x0000000000108000) 
//    12'h738 : LOC <=          63'b000000000000000000000000000000000000000001000001000000000000000; // D (0x0000000000208000) 
//    12'h74d : LOC <=          63'b000000000000000000000000000000000000000010000001000000000000000; // D (0x0000000000408000) 
//    12'h7a7 : LOC <=          63'b000000000000000000000000000000000000000100000001000000000000000; // D (0x0000000000808000) 
//    12'h673 : LOC <=          63'b000000000000000000000000000000000000001000000001000000000000000; // D (0x0000000001008000) 
//    12'h5db : LOC <=          63'b000000000000000000000000000000000000010000000001000000000000000; // D (0x0000000002008000) 
//    12'h28b : LOC <=          63'b000000000000000000000000000000000000100000000001000000000000000; // D (0x0000000004008000) 
//    12'hc2b : LOC <=          63'b000000000000000000000000000000000001000000000001000000000000000; // D (0x0000000008008000) 
//    12'h452 : LOC <=          63'b000000000000000000000000000000000010000000000001000000000000000; // D (0x0000000010008000) 
//    12'h199 : LOC <=          63'b000000000000000000000000000000000100000000000001000000000000000; // D (0x0000000020008000) 
//    12'ha0f : LOC <=          63'b000000000000000000000000000000001000000000000001000000000000000; // D (0x0000000040008000) 
//    12'h81a : LOC <=          63'b000000000000000000000000000000010000000000000001000000000000000; // D (0x0000000080008000) 
//    12'hc30 : LOC <=          63'b000000000000000000000000000000100000000000000001000000000000000; // D (0x0000000100008000) 
//    12'h464 : LOC <=          63'b000000000000000000000000000001000000000000000001000000000000000; // D (0x0000000200008000) 
//    12'h1f5 : LOC <=          63'b000000000000000000000000000010000000000000000001000000000000000; // D (0x0000000400008000) 
//    12'had7 : LOC <=          63'b000000000000000000000000000100000000000000000001000000000000000; // D (0x0000000800008000) 
//    12'h9aa : LOC <=          63'b000000000000000000000000001000000000000000000001000000000000000; // D (0x0000001000008000) 
//    12'hf50 : LOC <=          63'b000000000000000000000000010000000000000000000001000000000000000; // D (0x0000002000008000) 
//    12'h2a4 : LOC <=          63'b000000000000000000000000100000000000000000000001000000000000000; // D (0x0000004000008000) 
//    12'hc75 : LOC <=          63'b000000000000000000000001000000000000000000000001000000000000000; // D (0x0000008000008000) 
//    12'h4ee : LOC <=          63'b000000000000000000000010000000000000000000000001000000000000000; // D (0x0000010000008000) 
//    12'h0e1 : LOC <=          63'b000000000000000000000100000000000000000000000001000000000000000; // D (0x0000020000008000) 
//    12'h8ff : LOC <=          63'b000000000000000000001000000000000000000000000001000000000000000; // D (0x0000040000008000) 
//    12'hdfa : LOC <=          63'b000000000000000000010000000000000000000000000001000000000000000; // D (0x0000080000008000) 
//    12'h7f0 : LOC <=          63'b000000000000000000100000000000000000000000000001000000000000000; // D (0x0000100000008000) 
//    12'h6dd : LOC <=          63'b000000000000000001000000000000000000000000000001000000000000000; // D (0x0000200000008000) 
//    12'h487 : LOC <=          63'b000000000000000010000000000000000000000000000001000000000000000; // D (0x0000400000008000) 
//    12'h033 : LOC <=          63'b000000000000000100000000000000000000000000000001000000000000000; // D (0x0000800000008000) 
//    12'h95b : LOC <=          63'b000000000000001000000000000000000000000000000001000000000000000; // D (0x0001000000008000) 
//    12'heb2 : LOC <=          63'b000000000000010000000000000000000000000000000001000000000000000; // D (0x0002000000008000) 
//    12'h160 : LOC <=          63'b000000000000100000000000000000000000000000000001000000000000000; // D (0x0004000000008000) 
//    12'hbfd : LOC <=          63'b000000000001000000000000000000000000000000000001000000000000000; // D (0x0008000000008000) 
//    12'hbfe : LOC <=          63'b000000000010000000000000000000000000000000000001000000000000000; // D (0x0010000000008000) 
//    12'hbf8 : LOC <=          63'b000000000100000000000000000000000000000000000001000000000000000; // D (0x0020000000008000) 
//    12'hbf4 : LOC <=          63'b000000001000000000000000000000000000000000000001000000000000000; // D (0x0040000000008000) 
//    12'hbec : LOC <=          63'b000000010000000000000000000000000000000000000001000000000000000; // D (0x0080000000008000) 
//    12'hbdc : LOC <=          63'b000000100000000000000000000000000000000000000001000000000000000; // D (0x0100000000008000) 
//    12'hbbc : LOC <=          63'b000001000000000000000000000000000000000000000001000000000000000; // D (0x0200000000008000) 
//    12'hb7c : LOC <=          63'b000010000000000000000000000000000000000000000001000000000000000; // D (0x0400000000008000) 
//    12'hafc : LOC <=          63'b000100000000000000000000000000000000000000000001000000000000000; // D (0x0800000000008000) 
//    12'h9fc : LOC <=          63'b001000000000000000000000000000000000000000000001000000000000000; // D (0x1000000000008000) 
//    12'hffc : LOC <=          63'b010000000000000000000000000000000000000000000001000000000000000; // D (0x2000000000008000) 
//    12'h3fc : LOC <=          63'b100000000000000000000000000000000000000000000001000000000000000; // D (0x4000000000008000) 
    12'h7f8 : LOC <=          63'b000000000000000000000000000000000000000000000010000000000000001; // D (0x0000000000010001) 
    12'h8b3 : LOC <=          63'b000000000000000000000000000000000000000000000010000000000000010; // D (0x0000000000010002) 
    12'h31c : LOC <=          63'b000000000000000000000000000000000000000000000010000000000000100; // D (0x0000000000010004) 
    12'h17b : LOC <=          63'b000000000000000000000000000000000000000000000010000000000001000; // D (0x0000000000010008) 
    12'h5b5 : LOC <=          63'b000000000000000000000000000000000000000000000010000000000010000; // D (0x0000000000010010) 
    12'hc29 : LOC <=          63'b000000000000000000000000000000000000000000000010000000000100000; // D (0x0000000000010020) 
    12'ha28 : LOC <=          63'b000000000000000000000000000000000000000000000010000000001000000; // D (0x0000000000010040) 
    12'h62a : LOC <=          63'b000000000000000000000000000000000000000000000010000000010000000; // D (0x0000000000010080) 
    12'hb17 : LOC <=          63'b000000000000000000000000000000000000000000000010000000100000000; // D (0x0000000000010100) 
    12'h454 : LOC <=          63'b000000000000000000000000000000000000000000000010000001000000000; // D (0x0000000000010200) 
    12'hfeb : LOC <=          63'b000000000000000000000000000000000000000000000010000010000000000; // D (0x0000000000010400) 
    12'hdac : LOC <=          63'b000000000000000000000000000000000000000000000010000100000000000; // D (0x0000000000010800) 
    12'h922 : LOC <=          63'b000000000000000000000000000000000000000000000010001000000000000; // D (0x0000000000011000) 
    12'h03e : LOC <=          63'b000000000000000000000000000000000000000000000010010000000000000; // D (0x0000000000012000) 
    12'h73f : LOC <=          63'b000000000000000000000000000000000000000000000010100000000000000; // D (0x0000000000014000) 
    12'h93d : LOC <=          63'b000000000000000000000000000000000000000000000011000000000000000; // D (0x0000000000018000) 
    12'h2c1 : LOC <=          63'b000000000000000000000000000000000000000000000010000000000000000; // S (0x0000000000010000) 
//    12'h743 : LOC <=          63'b000000000000000000000000000000000000000000000110000000000000000; // D (0x0000000000030000) 
//    12'h9c5 : LOC <=          63'b000000000000000000000000000000000000000000001010000000000000000; // D (0x0000000000050000) 
//    12'h1f0 : LOC <=          63'b000000000000000000000000000000000000000000010010000000000000000; // D (0x0000000000090000) 
//    12'h4a3 : LOC <=          63'b000000000000000000000000000000000000000000100010000000000000000; // D (0x0000000000110000) 
//    12'he05 : LOC <=          63'b000000000000000000000000000000000000000001000010000000000000000; // D (0x0000000000210000) 
//    12'he70 : LOC <=          63'b000000000000000000000000000000000000000010000010000000000000000; // D (0x0000000000410000) 
//    12'he9a : LOC <=          63'b000000000000000000000000000000000000000100000010000000000000000; // D (0x0000000000810000) 
//    12'hf4e : LOC <=          63'b000000000000000000000000000000000000001000000010000000000000000; // D (0x0000000001010000) 
//    12'hce6 : LOC <=          63'b000000000000000000000000000000000000010000000010000000000000000; // D (0x0000000002010000) 
//    12'hbb6 : LOC <=          63'b000000000000000000000000000000000000100000000010000000000000000; // D (0x0000000004010000) 
//    12'h516 : LOC <=          63'b000000000000000000000000000000000001000000000010000000000000000; // D (0x0000000008010000) 
//    12'hd6f : LOC <=          63'b000000000000000000000000000000000010000000000010000000000000000; // D (0x0000000010010000) 
//    12'h8a4 : LOC <=          63'b000000000000000000000000000000000100000000000010000000000000000; // D (0x0000000020010000) 
//    12'h332 : LOC <=          63'b000000000000000000000000000000001000000000000010000000000000000; // D (0x0000000040010000) 
//    12'h127 : LOC <=          63'b000000000000000000000000000000010000000000000010000000000000000; // D (0x0000000080010000) 
//    12'h50d : LOC <=          63'b000000000000000000000000000000100000000000000010000000000000000; // D (0x0000000100010000) 
//    12'hd59 : LOC <=          63'b000000000000000000000000000001000000000000000010000000000000000; // D (0x0000000200010000) 
//    12'h8c8 : LOC <=          63'b000000000000000000000000000010000000000000000010000000000000000; // D (0x0000000400010000) 
//    12'h3ea : LOC <=          63'b000000000000000000000000000100000000000000000010000000000000000; // D (0x0000000800010000) 
//    12'h097 : LOC <=          63'b000000000000000000000000001000000000000000000010000000000000000; // D (0x0000001000010000) 
//    12'h66d : LOC <=          63'b000000000000000000000000010000000000000000000010000000000000000; // D (0x0000002000010000) 
//    12'hb99 : LOC <=          63'b000000000000000000000000100000000000000000000010000000000000000; // D (0x0000004000010000) 
//    12'h548 : LOC <=          63'b000000000000000000000001000000000000000000000010000000000000000; // D (0x0000008000010000) 
//    12'hdd3 : LOC <=          63'b000000000000000000000010000000000000000000000010000000000000000; // D (0x0000010000010000) 
//    12'h9dc : LOC <=          63'b000000000000000000000100000000000000000000000010000000000000000; // D (0x0000020000010000) 
//    12'h1c2 : LOC <=          63'b000000000000000000001000000000000000000000000010000000000000000; // D (0x0000040000010000) 
//    12'h4c7 : LOC <=          63'b000000000000000000010000000000000000000000000010000000000000000; // D (0x0000080000010000) 
//    12'hecd : LOC <=          63'b000000000000000000100000000000000000000000000010000000000000000; // D (0x0000100000010000) 
//    12'hfe0 : LOC <=          63'b000000000000000001000000000000000000000000000010000000000000000; // D (0x0000200000010000) 
//    12'hdba : LOC <=          63'b000000000000000010000000000000000000000000000010000000000000000; // D (0x0000400000010000) 
//    12'h90e : LOC <=          63'b000000000000000100000000000000000000000000000010000000000000000; // D (0x0000800000010000) 
//    12'h066 : LOC <=          63'b000000000000001000000000000000000000000000000010000000000000000; // D (0x0001000000010000) 
//    12'h78f : LOC <=          63'b000000000000010000000000000000000000000000000010000000000000000; // D (0x0002000000010000) 
//    12'h85d : LOC <=          63'b000000000000100000000000000000000000000000000010000000000000000; // D (0x0004000000010000) 
//    12'h2c0 : LOC <=          63'b000000000001000000000000000000000000000000000010000000000000000; // D (0x0008000000010000) 
//    12'h2c3 : LOC <=          63'b000000000010000000000000000000000000000000000010000000000000000; // D (0x0010000000010000) 
//    12'h2c5 : LOC <=          63'b000000000100000000000000000000000000000000000010000000000000000; // D (0x0020000000010000) 
//    12'h2c9 : LOC <=          63'b000000001000000000000000000000000000000000000010000000000000000; // D (0x0040000000010000) 
//    12'h2d1 : LOC <=          63'b000000010000000000000000000000000000000000000010000000000000000; // D (0x0080000000010000) 
//    12'h2e1 : LOC <=          63'b000000100000000000000000000000000000000000000010000000000000000; // D (0x0100000000010000) 
//    12'h281 : LOC <=          63'b000001000000000000000000000000000000000000000010000000000000000; // D (0x0200000000010000) 
//    12'h241 : LOC <=          63'b000010000000000000000000000000000000000000000010000000000000000; // D (0x0400000000010000) 
//    12'h3c1 : LOC <=          63'b000100000000000000000000000000000000000000000010000000000000000; // D (0x0800000000010000) 
//    12'h0c1 : LOC <=          63'b001000000000000000000000000000000000000000000010000000000000000; // D (0x1000000000010000) 
//    12'h6c1 : LOC <=          63'b010000000000000000000000000000000000000000000010000000000000000; // D (0x2000000000010000) 
//    12'hac1 : LOC <=          63'b100000000000000000000000000000000000000000000010000000000000000; // D (0x4000000000010000) 
    12'h0bb : LOC <=          63'b000000000000000000000000000000000000000000000100000000000000001; // D (0x0000000000020001) 
    12'hff0 : LOC <=          63'b000000000000000000000000000000000000000000000100000000000000010; // D (0x0000000000020002) 
    12'h45f : LOC <=          63'b000000000000000000000000000000000000000000000100000000000000100; // D (0x0000000000020004) 
    12'h638 : LOC <=          63'b000000000000000000000000000000000000000000000100000000000001000; // D (0x0000000000020008) 
    12'h2f6 : LOC <=          63'b000000000000000000000000000000000000000000000100000000000010000; // D (0x0000000000020010) 
    12'hb6a : LOC <=          63'b000000000000000000000000000000000000000000000100000000000100000; // D (0x0000000000020020) 
    12'hd6b : LOC <=          63'b000000000000000000000000000000000000000000000100000000001000000; // D (0x0000000000020040) 
    12'h169 : LOC <=          63'b000000000000000000000000000000000000000000000100000000010000000; // D (0x0000000000020080) 
    12'hc54 : LOC <=          63'b000000000000000000000000000000000000000000000100000000100000000; // D (0x0000000000020100) 
    12'h317 : LOC <=          63'b000000000000000000000000000000000000000000000100000001000000000; // D (0x0000000000020200) 
    12'h8a8 : LOC <=          63'b000000000000000000000000000000000000000000000100000010000000000; // D (0x0000000000020400) 
    12'haef : LOC <=          63'b000000000000000000000000000000000000000000000100000100000000000; // D (0x0000000000020800) 
    12'he61 : LOC <=          63'b000000000000000000000000000000000000000000000100001000000000000; // D (0x0000000000021000) 
    12'h77d : LOC <=          63'b000000000000000000000000000000000000000000000100010000000000000; // D (0x0000000000022000) 
    12'h07c : LOC <=          63'b000000000000000000000000000000000000000000000100100000000000000; // D (0x0000000000024000) 
    12'he7e : LOC <=          63'b000000000000000000000000000000000000000000000101000000000000000; // D (0x0000000000028000) 
    12'h743 : LOC <=          63'b000000000000000000000000000000000000000000000110000000000000000; // D (0x0000000000030000) 
    12'h582 : LOC <=          63'b000000000000000000000000000000000000000000000100000000000000000; // S (0x0000000000020000) 
//    12'he86 : LOC <=          63'b000000000000000000000000000000000000000000001100000000000000000; // D (0x0000000000060000) 
//    12'h6b3 : LOC <=          63'b000000000000000000000000000000000000000000010100000000000000000; // D (0x00000000000a0000) 
//    12'h3e0 : LOC <=          63'b000000000000000000000000000000000000000000100100000000000000000; // D (0x0000000000120000) 
//    12'h946 : LOC <=          63'b000000000000000000000000000000000000000001000100000000000000000; // D (0x0000000000220000) 
//    12'h933 : LOC <=          63'b000000000000000000000000000000000000000010000100000000000000000; // D (0x0000000000420000) 
//    12'h9d9 : LOC <=          63'b000000000000000000000000000000000000000100000100000000000000000; // D (0x0000000000820000) 
//    12'h80d : LOC <=          63'b000000000000000000000000000000000000001000000100000000000000000; // D (0x0000000001020000) 
//    12'hba5 : LOC <=          63'b000000000000000000000000000000000000010000000100000000000000000; // D (0x0000000002020000) 
//    12'hcf5 : LOC <=          63'b000000000000000000000000000000000000100000000100000000000000000; // D (0x0000000004020000) 
//    12'h255 : LOC <=          63'b000000000000000000000000000000000001000000000100000000000000000; // D (0x0000000008020000) 
//    12'ha2c : LOC <=          63'b000000000000000000000000000000000010000000000100000000000000000; // D (0x0000000010020000) 
//    12'hfe7 : LOC <=          63'b000000000000000000000000000000000100000000000100000000000000000; // D (0x0000000020020000) 
//    12'h471 : LOC <=          63'b000000000000000000000000000000001000000000000100000000000000000; // D (0x0000000040020000) 
//    12'h664 : LOC <=          63'b000000000000000000000000000000010000000000000100000000000000000; // D (0x0000000080020000) 
//    12'h24e : LOC <=          63'b000000000000000000000000000000100000000000000100000000000000000; // D (0x0000000100020000) 
//    12'ha1a : LOC <=          63'b000000000000000000000000000001000000000000000100000000000000000; // D (0x0000000200020000) 
//    12'hf8b : LOC <=          63'b000000000000000000000000000010000000000000000100000000000000000; // D (0x0000000400020000) 
//    12'h4a9 : LOC <=          63'b000000000000000000000000000100000000000000000100000000000000000; // D (0x0000000800020000) 
//    12'h7d4 : LOC <=          63'b000000000000000000000000001000000000000000000100000000000000000; // D (0x0000001000020000) 
//    12'h12e : LOC <=          63'b000000000000000000000000010000000000000000000100000000000000000; // D (0x0000002000020000) 
//    12'hcda : LOC <=          63'b000000000000000000000000100000000000000000000100000000000000000; // D (0x0000004000020000) 
//    12'h20b : LOC <=          63'b000000000000000000000001000000000000000000000100000000000000000; // D (0x0000008000020000) 
//    12'ha90 : LOC <=          63'b000000000000000000000010000000000000000000000100000000000000000; // D (0x0000010000020000) 
//    12'he9f : LOC <=          63'b000000000000000000000100000000000000000000000100000000000000000; // D (0x0000020000020000) 
//    12'h681 : LOC <=          63'b000000000000000000001000000000000000000000000100000000000000000; // D (0x0000040000020000) 
//    12'h384 : LOC <=          63'b000000000000000000010000000000000000000000000100000000000000000; // D (0x0000080000020000) 
//    12'h98e : LOC <=          63'b000000000000000000100000000000000000000000000100000000000000000; // D (0x0000100000020000) 
//    12'h8a3 : LOC <=          63'b000000000000000001000000000000000000000000000100000000000000000; // D (0x0000200000020000) 
//    12'haf9 : LOC <=          63'b000000000000000010000000000000000000000000000100000000000000000; // D (0x0000400000020000) 
//    12'he4d : LOC <=          63'b000000000000000100000000000000000000000000000100000000000000000; // D (0x0000800000020000) 
//    12'h725 : LOC <=          63'b000000000000001000000000000000000000000000000100000000000000000; // D (0x0001000000020000) 
//    12'h0cc : LOC <=          63'b000000000000010000000000000000000000000000000100000000000000000; // D (0x0002000000020000) 
//    12'hf1e : LOC <=          63'b000000000000100000000000000000000000000000000100000000000000000; // D (0x0004000000020000) 
//    12'h583 : LOC <=          63'b000000000001000000000000000000000000000000000100000000000000000; // D (0x0008000000020000) 
//    12'h580 : LOC <=          63'b000000000010000000000000000000000000000000000100000000000000000; // D (0x0010000000020000) 
//    12'h586 : LOC <=          63'b000000000100000000000000000000000000000000000100000000000000000; // D (0x0020000000020000) 
//    12'h58a : LOC <=          63'b000000001000000000000000000000000000000000000100000000000000000; // D (0x0040000000020000) 
//    12'h592 : LOC <=          63'b000000010000000000000000000000000000000000000100000000000000000; // D (0x0080000000020000) 
//    12'h5a2 : LOC <=          63'b000000100000000000000000000000000000000000000100000000000000000; // D (0x0100000000020000) 
//    12'h5c2 : LOC <=          63'b000001000000000000000000000000000000000000000100000000000000000; // D (0x0200000000020000) 
//    12'h502 : LOC <=          63'b000010000000000000000000000000000000000000000100000000000000000; // D (0x0400000000020000) 
//    12'h482 : LOC <=          63'b000100000000000000000000000000000000000000000100000000000000000; // D (0x0800000000020000) 
//    12'h782 : LOC <=          63'b001000000000000000000000000000000000000000000100000000000000000; // D (0x1000000000020000) 
//    12'h182 : LOC <=          63'b010000000000000000000000000000000000000000000100000000000000000; // D (0x2000000000020000) 
//    12'hd82 : LOC <=          63'b100000000000000000000000000000000000000000000100000000000000000; // D (0x4000000000020000) 
    12'he3d : LOC <=          63'b000000000000000000000000000000000000000000001000000000000000001; // D (0x0000000000040001) 
    12'h176 : LOC <=          63'b000000000000000000000000000000000000000000001000000000000000010; // D (0x0000000000040002) 
    12'had9 : LOC <=          63'b000000000000000000000000000000000000000000001000000000000000100; // D (0x0000000000040004) 
    12'h8be : LOC <=          63'b000000000000000000000000000000000000000000001000000000000001000; // D (0x0000000000040008) 
    12'hc70 : LOC <=          63'b000000000000000000000000000000000000000000001000000000000010000; // D (0x0000000000040010) 
    12'h5ec : LOC <=          63'b000000000000000000000000000000000000000000001000000000000100000; // D (0x0000000000040020) 
    12'h3ed : LOC <=          63'b000000000000000000000000000000000000000000001000000000001000000; // D (0x0000000000040040) 
    12'hfef : LOC <=          63'b000000000000000000000000000000000000000000001000000000010000000; // D (0x0000000000040080) 
    12'h2d2 : LOC <=          63'b000000000000000000000000000000000000000000001000000000100000000; // D (0x0000000000040100) 
    12'hd91 : LOC <=          63'b000000000000000000000000000000000000000000001000000001000000000; // D (0x0000000000040200) 
    12'h62e : LOC <=          63'b000000000000000000000000000000000000000000001000000010000000000; // D (0x0000000000040400) 
    12'h469 : LOC <=          63'b000000000000000000000000000000000000000000001000000100000000000; // D (0x0000000000040800) 
    12'h0e7 : LOC <=          63'b000000000000000000000000000000000000000000001000001000000000000; // D (0x0000000000041000) 
    12'h9fb : LOC <=          63'b000000000000000000000000000000000000000000001000010000000000000; // D (0x0000000000042000) 
    12'hefa : LOC <=          63'b000000000000000000000000000000000000000000001000100000000000000; // D (0x0000000000044000) 
    12'h0f8 : LOC <=          63'b000000000000000000000000000000000000000000001001000000000000000; // D (0x0000000000048000) 
    12'h9c5 : LOC <=          63'b000000000000000000000000000000000000000000001010000000000000000; // D (0x0000000000050000) 
    12'he86 : LOC <=          63'b000000000000000000000000000000000000000000001100000000000000000; // D (0x0000000000060000) 
    12'hb04 : LOC <=          63'b000000000000000000000000000000000000000000001000000000000000000; // S (0x0000000000040000) 
//    12'h835 : LOC <=          63'b000000000000000000000000000000000000000000011000000000000000000; // D (0x00000000000c0000) 
//    12'hd66 : LOC <=          63'b000000000000000000000000000000000000000000101000000000000000000; // D (0x0000000000140000) 
//    12'h7c0 : LOC <=          63'b000000000000000000000000000000000000000001001000000000000000000; // D (0x0000000000240000) 
//    12'h7b5 : LOC <=          63'b000000000000000000000000000000000000000010001000000000000000000; // D (0x0000000000440000) 
//    12'h75f : LOC <=          63'b000000000000000000000000000000000000000100001000000000000000000; // D (0x0000000000840000) 
//    12'h68b : LOC <=          63'b000000000000000000000000000000000000001000001000000000000000000; // D (0x0000000001040000) 
//    12'h523 : LOC <=          63'b000000000000000000000000000000000000010000001000000000000000000; // D (0x0000000002040000) 
//    12'h273 : LOC <=          63'b000000000000000000000000000000000000100000001000000000000000000; // D (0x0000000004040000) 
//    12'hcd3 : LOC <=          63'b000000000000000000000000000000000001000000001000000000000000000; // D (0x0000000008040000) 
//    12'h4aa : LOC <=          63'b000000000000000000000000000000000010000000001000000000000000000; // D (0x0000000010040000) 
//    12'h161 : LOC <=          63'b000000000000000000000000000000000100000000001000000000000000000; // D (0x0000000020040000) 
//    12'haf7 : LOC <=          63'b000000000000000000000000000000001000000000001000000000000000000; // D (0x0000000040040000) 
//    12'h8e2 : LOC <=          63'b000000000000000000000000000000010000000000001000000000000000000; // D (0x0000000080040000) 
//    12'hcc8 : LOC <=          63'b000000000000000000000000000000100000000000001000000000000000000; // D (0x0000000100040000) 
//    12'h49c : LOC <=          63'b000000000000000000000000000001000000000000001000000000000000000; // D (0x0000000200040000) 
//    12'h10d : LOC <=          63'b000000000000000000000000000010000000000000001000000000000000000; // D (0x0000000400040000) 
//    12'ha2f : LOC <=          63'b000000000000000000000000000100000000000000001000000000000000000; // D (0x0000000800040000) 
//    12'h952 : LOC <=          63'b000000000000000000000000001000000000000000001000000000000000000; // D (0x0000001000040000) 
//    12'hfa8 : LOC <=          63'b000000000000000000000000010000000000000000001000000000000000000; // D (0x0000002000040000) 
//    12'h25c : LOC <=          63'b000000000000000000000000100000000000000000001000000000000000000; // D (0x0000004000040000) 
//    12'hc8d : LOC <=          63'b000000000000000000000001000000000000000000001000000000000000000; // D (0x0000008000040000) 
//    12'h416 : LOC <=          63'b000000000000000000000010000000000000000000001000000000000000000; // D (0x0000010000040000) 
//    12'h019 : LOC <=          63'b000000000000000000000100000000000000000000001000000000000000000; // D (0x0000020000040000) 
//    12'h807 : LOC <=          63'b000000000000000000001000000000000000000000001000000000000000000; // D (0x0000040000040000) 
//    12'hd02 : LOC <=          63'b000000000000000000010000000000000000000000001000000000000000000; // D (0x0000080000040000) 
//    12'h708 : LOC <=          63'b000000000000000000100000000000000000000000001000000000000000000; // D (0x0000100000040000) 
//    12'h625 : LOC <=          63'b000000000000000001000000000000000000000000001000000000000000000; // D (0x0000200000040000) 
//    12'h47f : LOC <=          63'b000000000000000010000000000000000000000000001000000000000000000; // D (0x0000400000040000) 
//    12'h0cb : LOC <=          63'b000000000000000100000000000000000000000000001000000000000000000; // D (0x0000800000040000) 
//    12'h9a3 : LOC <=          63'b000000000000001000000000000000000000000000001000000000000000000; // D (0x0001000000040000) 
//    12'he4a : LOC <=          63'b000000000000010000000000000000000000000000001000000000000000000; // D (0x0002000000040000) 
//    12'h198 : LOC <=          63'b000000000000100000000000000000000000000000001000000000000000000; // D (0x0004000000040000) 
//    12'hb05 : LOC <=          63'b000000000001000000000000000000000000000000001000000000000000000; // D (0x0008000000040000) 
//    12'hb06 : LOC <=          63'b000000000010000000000000000000000000000000001000000000000000000; // D (0x0010000000040000) 
//    12'hb00 : LOC <=          63'b000000000100000000000000000000000000000000001000000000000000000; // D (0x0020000000040000) 
//    12'hb0c : LOC <=          63'b000000001000000000000000000000000000000000001000000000000000000; // D (0x0040000000040000) 
//    12'hb14 : LOC <=          63'b000000010000000000000000000000000000000000001000000000000000000; // D (0x0080000000040000) 
//    12'hb24 : LOC <=          63'b000000100000000000000000000000000000000000001000000000000000000; // D (0x0100000000040000) 
//    12'hb44 : LOC <=          63'b000001000000000000000000000000000000000000001000000000000000000; // D (0x0200000000040000) 
//    12'hb84 : LOC <=          63'b000010000000000000000000000000000000000000001000000000000000000; // D (0x0400000000040000) 
//    12'ha04 : LOC <=          63'b000100000000000000000000000000000000000000001000000000000000000; // D (0x0800000000040000) 
//    12'h904 : LOC <=          63'b001000000000000000000000000000000000000000001000000000000000000; // D (0x1000000000040000) 
//    12'hf04 : LOC <=          63'b010000000000000000000000000000000000000000001000000000000000000; // D (0x2000000000040000) 
//    12'h304 : LOC <=          63'b100000000000000000000000000000000000000000001000000000000000000; // D (0x4000000000040000) 
    12'h608 : LOC <=          63'b000000000000000000000000000000000000000000010000000000000000001; // D (0x0000000000080001) 
    12'h943 : LOC <=          63'b000000000000000000000000000000000000000000010000000000000000010; // D (0x0000000000080002) 
    12'h2ec : LOC <=          63'b000000000000000000000000000000000000000000010000000000000000100; // D (0x0000000000080004) 
    12'h08b : LOC <=          63'b000000000000000000000000000000000000000000010000000000000001000; // D (0x0000000000080008) 
    12'h445 : LOC <=          63'b000000000000000000000000000000000000000000010000000000000010000; // D (0x0000000000080010) 
    12'hdd9 : LOC <=          63'b000000000000000000000000000000000000000000010000000000000100000; // D (0x0000000000080020) 
    12'hbd8 : LOC <=          63'b000000000000000000000000000000000000000000010000000000001000000; // D (0x0000000000080040) 
    12'h7da : LOC <=          63'b000000000000000000000000000000000000000000010000000000010000000; // D (0x0000000000080080) 
    12'hae7 : LOC <=          63'b000000000000000000000000000000000000000000010000000000100000000; // D (0x0000000000080100) 
    12'h5a4 : LOC <=          63'b000000000000000000000000000000000000000000010000000001000000000; // D (0x0000000000080200) 
    12'he1b : LOC <=          63'b000000000000000000000000000000000000000000010000000010000000000; // D (0x0000000000080400) 
    12'hc5c : LOC <=          63'b000000000000000000000000000000000000000000010000000100000000000; // D (0x0000000000080800) 
    12'h8d2 : LOC <=          63'b000000000000000000000000000000000000000000010000001000000000000; // D (0x0000000000081000) 
    12'h1ce : LOC <=          63'b000000000000000000000000000000000000000000010000010000000000000; // D (0x0000000000082000) 
    12'h6cf : LOC <=          63'b000000000000000000000000000000000000000000010000100000000000000; // D (0x0000000000084000) 
    12'h8cd : LOC <=          63'b000000000000000000000000000000000000000000010001000000000000000; // D (0x0000000000088000) 
    12'h1f0 : LOC <=          63'b000000000000000000000000000000000000000000010010000000000000000; // D (0x0000000000090000) 
    12'h6b3 : LOC <=          63'b000000000000000000000000000000000000000000010100000000000000000; // D (0x00000000000a0000) 
    12'h835 : LOC <=          63'b000000000000000000000000000000000000000000011000000000000000000; // D (0x00000000000c0000) 
    12'h331 : LOC <=          63'b000000000000000000000000000000000000000000010000000000000000000; // S (0x0000000000080000) 
//    12'h553 : LOC <=          63'b000000000000000000000000000000000000000000110000000000000000000; // D (0x0000000000180000) 
//    12'hff5 : LOC <=          63'b000000000000000000000000000000000000000001010000000000000000000; // D (0x0000000000280000) 
//    12'hf80 : LOC <=          63'b000000000000000000000000000000000000000010010000000000000000000; // D (0x0000000000480000) 
//    12'hf6a : LOC <=          63'b000000000000000000000000000000000000000100010000000000000000000; // D (0x0000000000880000) 
//    12'hebe : LOC <=          63'b000000000000000000000000000000000000001000010000000000000000000; // D (0x0000000001080000) 
//    12'hd16 : LOC <=          63'b000000000000000000000000000000000000010000010000000000000000000; // D (0x0000000002080000) 
//    12'ha46 : LOC <=          63'b000000000000000000000000000000000000100000010000000000000000000; // D (0x0000000004080000) 
//    12'h4e6 : LOC <=          63'b000000000000000000000000000000000001000000010000000000000000000; // D (0x0000000008080000) 
//    12'hc9f : LOC <=          63'b000000000000000000000000000000000010000000010000000000000000000; // D (0x0000000010080000) 
//    12'h954 : LOC <=          63'b000000000000000000000000000000000100000000010000000000000000000; // D (0x0000000020080000) 
//    12'h2c2 : LOC <=          63'b000000000000000000000000000000001000000000010000000000000000000; // D (0x0000000040080000) 
//    12'h0d7 : LOC <=          63'b000000000000000000000000000000010000000000010000000000000000000; // D (0x0000000080080000) 
//    12'h4fd : LOC <=          63'b000000000000000000000000000000100000000000010000000000000000000; // D (0x0000000100080000) 
//    12'hca9 : LOC <=          63'b000000000000000000000000000001000000000000010000000000000000000; // D (0x0000000200080000) 
//    12'h938 : LOC <=          63'b000000000000000000000000000010000000000000010000000000000000000; // D (0x0000000400080000) 
//    12'h21a : LOC <=          63'b000000000000000000000000000100000000000000010000000000000000000; // D (0x0000000800080000) 
//    12'h167 : LOC <=          63'b000000000000000000000000001000000000000000010000000000000000000; // D (0x0000001000080000) 
//    12'h79d : LOC <=          63'b000000000000000000000000010000000000000000010000000000000000000; // D (0x0000002000080000) 
//    12'ha69 : LOC <=          63'b000000000000000000000000100000000000000000010000000000000000000; // D (0x0000004000080000) 
//    12'h4b8 : LOC <=          63'b000000000000000000000001000000000000000000010000000000000000000; // D (0x0000008000080000) 
//    12'hc23 : LOC <=          63'b000000000000000000000010000000000000000000010000000000000000000; // D (0x0000010000080000) 
//    12'h82c : LOC <=          63'b000000000000000000000100000000000000000000010000000000000000000; // D (0x0000020000080000) 
//    12'h032 : LOC <=          63'b000000000000000000001000000000000000000000010000000000000000000; // D (0x0000040000080000) 
//    12'h537 : LOC <=          63'b000000000000000000010000000000000000000000010000000000000000000; // D (0x0000080000080000) 
//    12'hf3d : LOC <=          63'b000000000000000000100000000000000000000000010000000000000000000; // D (0x0000100000080000) 
//    12'he10 : LOC <=          63'b000000000000000001000000000000000000000000010000000000000000000; // D (0x0000200000080000) 
//    12'hc4a : LOC <=          63'b000000000000000010000000000000000000000000010000000000000000000; // D (0x0000400000080000) 
//    12'h8fe : LOC <=          63'b000000000000000100000000000000000000000000010000000000000000000; // D (0x0000800000080000) 
//    12'h196 : LOC <=          63'b000000000000001000000000000000000000000000010000000000000000000; // D (0x0001000000080000) 
//    12'h67f : LOC <=          63'b000000000000010000000000000000000000000000010000000000000000000; // D (0x0002000000080000) 
//    12'h9ad : LOC <=          63'b000000000000100000000000000000000000000000010000000000000000000; // D (0x0004000000080000) 
//    12'h330 : LOC <=          63'b000000000001000000000000000000000000000000010000000000000000000; // D (0x0008000000080000) 
//    12'h333 : LOC <=          63'b000000000010000000000000000000000000000000010000000000000000000; // D (0x0010000000080000) 
//    12'h335 : LOC <=          63'b000000000100000000000000000000000000000000010000000000000000000; // D (0x0020000000080000) 
//    12'h339 : LOC <=          63'b000000001000000000000000000000000000000000010000000000000000000; // D (0x0040000000080000) 
//    12'h321 : LOC <=          63'b000000010000000000000000000000000000000000010000000000000000000; // D (0x0080000000080000) 
//    12'h311 : LOC <=          63'b000000100000000000000000000000000000000000010000000000000000000; // D (0x0100000000080000) 
//    12'h371 : LOC <=          63'b000001000000000000000000000000000000000000010000000000000000000; // D (0x0200000000080000) 
//    12'h3b1 : LOC <=          63'b000010000000000000000000000000000000000000010000000000000000000; // D (0x0400000000080000) 
//    12'h231 : LOC <=          63'b000100000000000000000000000000000000000000010000000000000000000; // D (0x0800000000080000) 
//    12'h131 : LOC <=          63'b001000000000000000000000000000000000000000010000000000000000000; // D (0x1000000000080000) 
//    12'h731 : LOC <=          63'b010000000000000000000000000000000000000000010000000000000000000; // D (0x2000000000080000) 
//    12'hb31 : LOC <=          63'b100000000000000000000000000000000000000000010000000000000000000; // D (0x4000000000080000) 
    12'h35b : LOC <=          63'b000000000000000000000000000000000000000000100000000000000000001; // D (0x0000000000100001) 
    12'hc10 : LOC <=          63'b000000000000000000000000000000000000000000100000000000000000010; // D (0x0000000000100002) 
    12'h7bf : LOC <=          63'b000000000000000000000000000000000000000000100000000000000000100; // D (0x0000000000100004) 
    12'h5d8 : LOC <=          63'b000000000000000000000000000000000000000000100000000000000001000; // D (0x0000000000100008) 
    12'h116 : LOC <=          63'b000000000000000000000000000000000000000000100000000000000010000; // D (0x0000000000100010) 
    12'h88a : LOC <=          63'b000000000000000000000000000000000000000000100000000000000100000; // D (0x0000000000100020) 
    12'he8b : LOC <=          63'b000000000000000000000000000000000000000000100000000000001000000; // D (0x0000000000100040) 
    12'h289 : LOC <=          63'b000000000000000000000000000000000000000000100000000000010000000; // D (0x0000000000100080) 
    12'hfb4 : LOC <=          63'b000000000000000000000000000000000000000000100000000000100000000; // D (0x0000000000100100) 
    12'h0f7 : LOC <=          63'b000000000000000000000000000000000000000000100000000001000000000; // D (0x0000000000100200) 
    12'hb48 : LOC <=          63'b000000000000000000000000000000000000000000100000000010000000000; // D (0x0000000000100400) 
    12'h90f : LOC <=          63'b000000000000000000000000000000000000000000100000000100000000000; // D (0x0000000000100800) 
    12'hd81 : LOC <=          63'b000000000000000000000000000000000000000000100000001000000000000; // D (0x0000000000101000) 
    12'h49d : LOC <=          63'b000000000000000000000000000000000000000000100000010000000000000; // D (0x0000000000102000) 
    12'h39c : LOC <=          63'b000000000000000000000000000000000000000000100000100000000000000; // D (0x0000000000104000) 
    12'hd9e : LOC <=          63'b000000000000000000000000000000000000000000100001000000000000000; // D (0x0000000000108000) 
    12'h4a3 : LOC <=          63'b000000000000000000000000000000000000000000100010000000000000000; // D (0x0000000000110000) 
    12'h3e0 : LOC <=          63'b000000000000000000000000000000000000000000100100000000000000000; // D (0x0000000000120000) 
    12'hd66 : LOC <=          63'b000000000000000000000000000000000000000000101000000000000000000; // D (0x0000000000140000) 
    12'h553 : LOC <=          63'b000000000000000000000000000000000000000000110000000000000000000; // D (0x0000000000180000) 
    12'h662 : LOC <=          63'b000000000000000000000000000000000000000000100000000000000000000; // S (0x0000000000100000) 
//    12'haa6 : LOC <=          63'b000000000000000000000000000000000000000001100000000000000000000; // D (0x0000000000300000) 
//    12'had3 : LOC <=          63'b000000000000000000000000000000000000000010100000000000000000000; // D (0x0000000000500000) 
//    12'ha39 : LOC <=          63'b000000000000000000000000000000000000000100100000000000000000000; // D (0x0000000000900000) 
//    12'hbed : LOC <=          63'b000000000000000000000000000000000000001000100000000000000000000; // D (0x0000000001100000) 
//    12'h845 : LOC <=          63'b000000000000000000000000000000000000010000100000000000000000000; // D (0x0000000002100000) 
//    12'hf15 : LOC <=          63'b000000000000000000000000000000000000100000100000000000000000000; // D (0x0000000004100000) 
//    12'h1b5 : LOC <=          63'b000000000000000000000000000000000001000000100000000000000000000; // D (0x0000000008100000) 
//    12'h9cc : LOC <=          63'b000000000000000000000000000000000010000000100000000000000000000; // D (0x0000000010100000) 
//    12'hc07 : LOC <=          63'b000000000000000000000000000000000100000000100000000000000000000; // D (0x0000000020100000) 
//    12'h791 : LOC <=          63'b000000000000000000000000000000001000000000100000000000000000000; // D (0x0000000040100000) 
//    12'h584 : LOC <=          63'b000000000000000000000000000000010000000000100000000000000000000; // D (0x0000000080100000) 
//    12'h1ae : LOC <=          63'b000000000000000000000000000000100000000000100000000000000000000; // D (0x0000000100100000) 
//    12'h9fa : LOC <=          63'b000000000000000000000000000001000000000000100000000000000000000; // D (0x0000000200100000) 
//    12'hc6b : LOC <=          63'b000000000000000000000000000010000000000000100000000000000000000; // D (0x0000000400100000) 
//    12'h749 : LOC <=          63'b000000000000000000000000000100000000000000100000000000000000000; // D (0x0000000800100000) 
//    12'h434 : LOC <=          63'b000000000000000000000000001000000000000000100000000000000000000; // D (0x0000001000100000) 
//    12'h2ce : LOC <=          63'b000000000000000000000000010000000000000000100000000000000000000; // D (0x0000002000100000) 
//    12'hf3a : LOC <=          63'b000000000000000000000000100000000000000000100000000000000000000; // D (0x0000004000100000) 
//    12'h1eb : LOC <=          63'b000000000000000000000001000000000000000000100000000000000000000; // D (0x0000008000100000) 
//    12'h970 : LOC <=          63'b000000000000000000000010000000000000000000100000000000000000000; // D (0x0000010000100000) 
//    12'hd7f : LOC <=          63'b000000000000000000000100000000000000000000100000000000000000000; // D (0x0000020000100000) 
//    12'h561 : LOC <=          63'b000000000000000000001000000000000000000000100000000000000000000; // D (0x0000040000100000) 
//    12'h064 : LOC <=          63'b000000000000000000010000000000000000000000100000000000000000000; // D (0x0000080000100000) 
//    12'ha6e : LOC <=          63'b000000000000000000100000000000000000000000100000000000000000000; // D (0x0000100000100000) 
//    12'hb43 : LOC <=          63'b000000000000000001000000000000000000000000100000000000000000000; // D (0x0000200000100000) 
//    12'h919 : LOC <=          63'b000000000000000010000000000000000000000000100000000000000000000; // D (0x0000400000100000) 
//    12'hdad : LOC <=          63'b000000000000000100000000000000000000000000100000000000000000000; // D (0x0000800000100000) 
//    12'h4c5 : LOC <=          63'b000000000000001000000000000000000000000000100000000000000000000; // D (0x0001000000100000) 
//    12'h32c : LOC <=          63'b000000000000010000000000000000000000000000100000000000000000000; // D (0x0002000000100000) 
//    12'hcfe : LOC <=          63'b000000000000100000000000000000000000000000100000000000000000000; // D (0x0004000000100000) 
//    12'h663 : LOC <=          63'b000000000001000000000000000000000000000000100000000000000000000; // D (0x0008000000100000) 
//    12'h660 : LOC <=          63'b000000000010000000000000000000000000000000100000000000000000000; // D (0x0010000000100000) 
//    12'h666 : LOC <=          63'b000000000100000000000000000000000000000000100000000000000000000; // D (0x0020000000100000) 
//    12'h66a : LOC <=          63'b000000001000000000000000000000000000000000100000000000000000000; // D (0x0040000000100000) 
//    12'h672 : LOC <=          63'b000000010000000000000000000000000000000000100000000000000000000; // D (0x0080000000100000) 
//    12'h642 : LOC <=          63'b000000100000000000000000000000000000000000100000000000000000000; // D (0x0100000000100000) 
//    12'h622 : LOC <=          63'b000001000000000000000000000000000000000000100000000000000000000; // D (0x0200000000100000) 
//    12'h6e2 : LOC <=          63'b000010000000000000000000000000000000000000100000000000000000000; // D (0x0400000000100000) 
//    12'h762 : LOC <=          63'b000100000000000000000000000000000000000000100000000000000000000; // D (0x0800000000100000) 
//    12'h462 : LOC <=          63'b001000000000000000000000000000000000000000100000000000000000000; // D (0x1000000000100000) 
//    12'h262 : LOC <=          63'b010000000000000000000000000000000000000000100000000000000000000; // D (0x2000000000100000) 
//    12'he62 : LOC <=          63'b100000000000000000000000000000000000000000100000000000000000000; // D (0x4000000000100000) 
    12'h9fd : LOC <=          63'b000000000000000000000000000000000000000001000000000000000000001; // D (0x0000000000200001) 
    12'h6b6 : LOC <=          63'b000000000000000000000000000000000000000001000000000000000000010; // D (0x0000000000200002) 
    12'hd19 : LOC <=          63'b000000000000000000000000000000000000000001000000000000000000100; // D (0x0000000000200004) 
    12'hf7e : LOC <=          63'b000000000000000000000000000000000000000001000000000000000001000; // D (0x0000000000200008) 
    12'hbb0 : LOC <=          63'b000000000000000000000000000000000000000001000000000000000010000; // D (0x0000000000200010) 
    12'h22c : LOC <=          63'b000000000000000000000000000000000000000001000000000000000100000; // D (0x0000000000200020) 
    12'h42d : LOC <=          63'b000000000000000000000000000000000000000001000000000000001000000; // D (0x0000000000200040) 
    12'h82f : LOC <=          63'b000000000000000000000000000000000000000001000000000000010000000; // D (0x0000000000200080) 
    12'h512 : LOC <=          63'b000000000000000000000000000000000000000001000000000000100000000; // D (0x0000000000200100) 
    12'ha51 : LOC <=          63'b000000000000000000000000000000000000000001000000000001000000000; // D (0x0000000000200200) 
    12'h1ee : LOC <=          63'b000000000000000000000000000000000000000001000000000010000000000; // D (0x0000000000200400) 
    12'h3a9 : LOC <=          63'b000000000000000000000000000000000000000001000000000100000000000; // D (0x0000000000200800) 
    12'h727 : LOC <=          63'b000000000000000000000000000000000000000001000000001000000000000; // D (0x0000000000201000) 
    12'he3b : LOC <=          63'b000000000000000000000000000000000000000001000000010000000000000; // D (0x0000000000202000) 
    12'h93a : LOC <=          63'b000000000000000000000000000000000000000001000000100000000000000; // D (0x0000000000204000) 
    12'h738 : LOC <=          63'b000000000000000000000000000000000000000001000001000000000000000; // D (0x0000000000208000) 
    12'he05 : LOC <=          63'b000000000000000000000000000000000000000001000010000000000000000; // D (0x0000000000210000) 
    12'h946 : LOC <=          63'b000000000000000000000000000000000000000001000100000000000000000; // D (0x0000000000220000) 
    12'h7c0 : LOC <=          63'b000000000000000000000000000000000000000001001000000000000000000; // D (0x0000000000240000) 
    12'hff5 : LOC <=          63'b000000000000000000000000000000000000000001010000000000000000000; // D (0x0000000000280000) 
    12'haa6 : LOC <=          63'b000000000000000000000000000000000000000001100000000000000000000; // D (0x0000000000300000) 
    12'hcc4 : LOC <=          63'b000000000000000000000000000000000000000001000000000000000000000; // S (0x0000000000200000) 
//    12'h075 : LOC <=          63'b000000000000000000000000000000000000000011000000000000000000000; // D (0x0000000000600000) 
//    12'h09f : LOC <=          63'b000000000000000000000000000000000000000101000000000000000000000; // D (0x0000000000a00000) 
//    12'h14b : LOC <=          63'b000000000000000000000000000000000000001001000000000000000000000; // D (0x0000000001200000) 
//    12'h2e3 : LOC <=          63'b000000000000000000000000000000000000010001000000000000000000000; // D (0x0000000002200000) 
//    12'h5b3 : LOC <=          63'b000000000000000000000000000000000000100001000000000000000000000; // D (0x0000000004200000) 
//    12'hb13 : LOC <=          63'b000000000000000000000000000000000001000001000000000000000000000; // D (0x0000000008200000) 
//    12'h36a : LOC <=          63'b000000000000000000000000000000000010000001000000000000000000000; // D (0x0000000010200000) 
//    12'h6a1 : LOC <=          63'b000000000000000000000000000000000100000001000000000000000000000; // D (0x0000000020200000) 
//    12'hd37 : LOC <=          63'b000000000000000000000000000000001000000001000000000000000000000; // D (0x0000000040200000) 
//    12'hf22 : LOC <=          63'b000000000000000000000000000000010000000001000000000000000000000; // D (0x0000000080200000) 
//    12'hb08 : LOC <=          63'b000000000000000000000000000000100000000001000000000000000000000; // D (0x0000000100200000) 
//    12'h35c : LOC <=          63'b000000000000000000000000000001000000000001000000000000000000000; // D (0x0000000200200000) 
//    12'h6cd : LOC <=          63'b000000000000000000000000000010000000000001000000000000000000000; // D (0x0000000400200000) 
//    12'hdef : LOC <=          63'b000000000000000000000000000100000000000001000000000000000000000; // D (0x0000000800200000) 
//    12'he92 : LOC <=          63'b000000000000000000000000001000000000000001000000000000000000000; // D (0x0000001000200000) 
//    12'h868 : LOC <=          63'b000000000000000000000000010000000000000001000000000000000000000; // D (0x0000002000200000) 
//    12'h59c : LOC <=          63'b000000000000000000000000100000000000000001000000000000000000000; // D (0x0000004000200000) 
//    12'hb4d : LOC <=          63'b000000000000000000000001000000000000000001000000000000000000000; // D (0x0000008000200000) 
//    12'h3d6 : LOC <=          63'b000000000000000000000010000000000000000001000000000000000000000; // D (0x0000010000200000) 
//    12'h7d9 : LOC <=          63'b000000000000000000000100000000000000000001000000000000000000000; // D (0x0000020000200000) 
//    12'hfc7 : LOC <=          63'b000000000000000000001000000000000000000001000000000000000000000; // D (0x0000040000200000) 
//    12'hac2 : LOC <=          63'b000000000000000000010000000000000000000001000000000000000000000; // D (0x0000080000200000) 
//    12'h0c8 : LOC <=          63'b000000000000000000100000000000000000000001000000000000000000000; // D (0x0000100000200000) 
//    12'h1e5 : LOC <=          63'b000000000000000001000000000000000000000001000000000000000000000; // D (0x0000200000200000) 
//    12'h3bf : LOC <=          63'b000000000000000010000000000000000000000001000000000000000000000; // D (0x0000400000200000) 
//    12'h70b : LOC <=          63'b000000000000000100000000000000000000000001000000000000000000000; // D (0x0000800000200000) 
//    12'he63 : LOC <=          63'b000000000000001000000000000000000000000001000000000000000000000; // D (0x0001000000200000) 
//    12'h98a : LOC <=          63'b000000000000010000000000000000000000000001000000000000000000000; // D (0x0002000000200000) 
//    12'h658 : LOC <=          63'b000000000000100000000000000000000000000001000000000000000000000; // D (0x0004000000200000) 
//    12'hcc5 : LOC <=          63'b000000000001000000000000000000000000000001000000000000000000000; // D (0x0008000000200000) 
//    12'hcc6 : LOC <=          63'b000000000010000000000000000000000000000001000000000000000000000; // D (0x0010000000200000) 
//    12'hcc0 : LOC <=          63'b000000000100000000000000000000000000000001000000000000000000000; // D (0x0020000000200000) 
//    12'hccc : LOC <=          63'b000000001000000000000000000000000000000001000000000000000000000; // D (0x0040000000200000) 
//    12'hcd4 : LOC <=          63'b000000010000000000000000000000000000000001000000000000000000000; // D (0x0080000000200000) 
//    12'hce4 : LOC <=          63'b000000100000000000000000000000000000000001000000000000000000000; // D (0x0100000000200000) 
//    12'hc84 : LOC <=          63'b000001000000000000000000000000000000000001000000000000000000000; // D (0x0200000000200000) 
//    12'hc44 : LOC <=          63'b000010000000000000000000000000000000000001000000000000000000000; // D (0x0400000000200000) 
//    12'hdc4 : LOC <=          63'b000100000000000000000000000000000000000001000000000000000000000; // D (0x0800000000200000) 
//    12'hec4 : LOC <=          63'b001000000000000000000000000000000000000001000000000000000000000; // D (0x1000000000200000) 
//    12'h8c4 : LOC <=          63'b010000000000000000000000000000000000000001000000000000000000000; // D (0x2000000000200000) 
//    12'h4c4 : LOC <=          63'b100000000000000000000000000000000000000001000000000000000000000; // D (0x4000000000200000) 
    12'h988 : LOC <=          63'b000000000000000000000000000000000000000010000000000000000000001; // D (0x0000000000400001) 
    12'h6c3 : LOC <=          63'b000000000000000000000000000000000000000010000000000000000000010; // D (0x0000000000400002) 
    12'hd6c : LOC <=          63'b000000000000000000000000000000000000000010000000000000000000100; // D (0x0000000000400004) 
    12'hf0b : LOC <=          63'b000000000000000000000000000000000000000010000000000000000001000; // D (0x0000000000400008) 
    12'hbc5 : LOC <=          63'b000000000000000000000000000000000000000010000000000000000010000; // D (0x0000000000400010) 
    12'h259 : LOC <=          63'b000000000000000000000000000000000000000010000000000000000100000; // D (0x0000000000400020) 
    12'h458 : LOC <=          63'b000000000000000000000000000000000000000010000000000000001000000; // D (0x0000000000400040) 
    12'h85a : LOC <=          63'b000000000000000000000000000000000000000010000000000000010000000; // D (0x0000000000400080) 
    12'h567 : LOC <=          63'b000000000000000000000000000000000000000010000000000000100000000; // D (0x0000000000400100) 
    12'ha24 : LOC <=          63'b000000000000000000000000000000000000000010000000000001000000000; // D (0x0000000000400200) 
    12'h19b : LOC <=          63'b000000000000000000000000000000000000000010000000000010000000000; // D (0x0000000000400400) 
    12'h3dc : LOC <=          63'b000000000000000000000000000000000000000010000000000100000000000; // D (0x0000000000400800) 
    12'h752 : LOC <=          63'b000000000000000000000000000000000000000010000000001000000000000; // D (0x0000000000401000) 
    12'he4e : LOC <=          63'b000000000000000000000000000000000000000010000000010000000000000; // D (0x0000000000402000) 
    12'h94f : LOC <=          63'b000000000000000000000000000000000000000010000000100000000000000; // D (0x0000000000404000) 
    12'h74d : LOC <=          63'b000000000000000000000000000000000000000010000001000000000000000; // D (0x0000000000408000) 
    12'he70 : LOC <=          63'b000000000000000000000000000000000000000010000010000000000000000; // D (0x0000000000410000) 
    12'h933 : LOC <=          63'b000000000000000000000000000000000000000010000100000000000000000; // D (0x0000000000420000) 
    12'h7b5 : LOC <=          63'b000000000000000000000000000000000000000010001000000000000000000; // D (0x0000000000440000) 
    12'hf80 : LOC <=          63'b000000000000000000000000000000000000000010010000000000000000000; // D (0x0000000000480000) 
    12'had3 : LOC <=          63'b000000000000000000000000000000000000000010100000000000000000000; // D (0x0000000000500000) 
    12'h075 : LOC <=          63'b000000000000000000000000000000000000000011000000000000000000000; // D (0x0000000000600000) 
    12'hcb1 : LOC <=          63'b000000000000000000000000000000000000000010000000000000000000000; // S (0x0000000000400000) 
//    12'h0ea : LOC <=          63'b000000000000000000000000000000000000000110000000000000000000000; // D (0x0000000000c00000) 
//    12'h13e : LOC <=          63'b000000000000000000000000000000000000001010000000000000000000000; // D (0x0000000001400000) 
//    12'h296 : LOC <=          63'b000000000000000000000000000000000000010010000000000000000000000; // D (0x0000000002400000) 
//    12'h5c6 : LOC <=          63'b000000000000000000000000000000000000100010000000000000000000000; // D (0x0000000004400000) 
//    12'hb66 : LOC <=          63'b000000000000000000000000000000000001000010000000000000000000000; // D (0x0000000008400000) 
//    12'h31f : LOC <=          63'b000000000000000000000000000000000010000010000000000000000000000; // D (0x0000000010400000) 
//    12'h6d4 : LOC <=          63'b000000000000000000000000000000000100000010000000000000000000000; // D (0x0000000020400000) 
//    12'hd42 : LOC <=          63'b000000000000000000000000000000001000000010000000000000000000000; // D (0x0000000040400000) 
//    12'hf57 : LOC <=          63'b000000000000000000000000000000010000000010000000000000000000000; // D (0x0000000080400000) 
//    12'hb7d : LOC <=          63'b000000000000000000000000000000100000000010000000000000000000000; // D (0x0000000100400000) 
//    12'h329 : LOC <=          63'b000000000000000000000000000001000000000010000000000000000000000; // D (0x0000000200400000) 
//    12'h6b8 : LOC <=          63'b000000000000000000000000000010000000000010000000000000000000000; // D (0x0000000400400000) 
//    12'hd9a : LOC <=          63'b000000000000000000000000000100000000000010000000000000000000000; // D (0x0000000800400000) 
//    12'hee7 : LOC <=          63'b000000000000000000000000001000000000000010000000000000000000000; // D (0x0000001000400000) 
//    12'h81d : LOC <=          63'b000000000000000000000000010000000000000010000000000000000000000; // D (0x0000002000400000) 
//    12'h5e9 : LOC <=          63'b000000000000000000000000100000000000000010000000000000000000000; // D (0x0000004000400000) 
//    12'hb38 : LOC <=          63'b000000000000000000000001000000000000000010000000000000000000000; // D (0x0000008000400000) 
//    12'h3a3 : LOC <=          63'b000000000000000000000010000000000000000010000000000000000000000; // D (0x0000010000400000) 
//    12'h7ac : LOC <=          63'b000000000000000000000100000000000000000010000000000000000000000; // D (0x0000020000400000) 
//    12'hfb2 : LOC <=          63'b000000000000000000001000000000000000000010000000000000000000000; // D (0x0000040000400000) 
//    12'hab7 : LOC <=          63'b000000000000000000010000000000000000000010000000000000000000000; // D (0x0000080000400000) 
//    12'h0bd : LOC <=          63'b000000000000000000100000000000000000000010000000000000000000000; // D (0x0000100000400000) 
//    12'h190 : LOC <=          63'b000000000000000001000000000000000000000010000000000000000000000; // D (0x0000200000400000) 
//    12'h3ca : LOC <=          63'b000000000000000010000000000000000000000010000000000000000000000; // D (0x0000400000400000) 
//    12'h77e : LOC <=          63'b000000000000000100000000000000000000000010000000000000000000000; // D (0x0000800000400000) 
//    12'he16 : LOC <=          63'b000000000000001000000000000000000000000010000000000000000000000; // D (0x0001000000400000) 
//    12'h9ff : LOC <=          63'b000000000000010000000000000000000000000010000000000000000000000; // D (0x0002000000400000) 
//    12'h62d : LOC <=          63'b000000000000100000000000000000000000000010000000000000000000000; // D (0x0004000000400000) 
//    12'hcb0 : LOC <=          63'b000000000001000000000000000000000000000010000000000000000000000; // D (0x0008000000400000) 
//    12'hcb3 : LOC <=          63'b000000000010000000000000000000000000000010000000000000000000000; // D (0x0010000000400000) 
//    12'hcb5 : LOC <=          63'b000000000100000000000000000000000000000010000000000000000000000; // D (0x0020000000400000) 
//    12'hcb9 : LOC <=          63'b000000001000000000000000000000000000000010000000000000000000000; // D (0x0040000000400000) 
//    12'hca1 : LOC <=          63'b000000010000000000000000000000000000000010000000000000000000000; // D (0x0080000000400000) 
//    12'hc91 : LOC <=          63'b000000100000000000000000000000000000000010000000000000000000000; // D (0x0100000000400000) 
//    12'hcf1 : LOC <=          63'b000001000000000000000000000000000000000010000000000000000000000; // D (0x0200000000400000) 
//    12'hc31 : LOC <=          63'b000010000000000000000000000000000000000010000000000000000000000; // D (0x0400000000400000) 
//    12'hdb1 : LOC <=          63'b000100000000000000000000000000000000000010000000000000000000000; // D (0x0800000000400000) 
//    12'heb1 : LOC <=          63'b001000000000000000000000000000000000000010000000000000000000000; // D (0x1000000000400000) 
//    12'h8b1 : LOC <=          63'b010000000000000000000000000000000000000010000000000000000000000; // D (0x2000000000400000) 
//    12'h4b1 : LOC <=          63'b100000000000000000000000000000000000000010000000000000000000000; // D (0x4000000000400000) 
    12'h962 : LOC <=          63'b000000000000000000000000000000000000000100000000000000000000001; // D (0x0000000000800001) 
    12'h629 : LOC <=          63'b000000000000000000000000000000000000000100000000000000000000010; // D (0x0000000000800002) 
    12'hd86 : LOC <=          63'b000000000000000000000000000000000000000100000000000000000000100; // D (0x0000000000800004) 
    12'hfe1 : LOC <=          63'b000000000000000000000000000000000000000100000000000000000001000; // D (0x0000000000800008) 
    12'hb2f : LOC <=          63'b000000000000000000000000000000000000000100000000000000000010000; // D (0x0000000000800010) 
    12'h2b3 : LOC <=          63'b000000000000000000000000000000000000000100000000000000000100000; // D (0x0000000000800020) 
    12'h4b2 : LOC <=          63'b000000000000000000000000000000000000000100000000000000001000000; // D (0x0000000000800040) 
    12'h8b0 : LOC <=          63'b000000000000000000000000000000000000000100000000000000010000000; // D (0x0000000000800080) 
    12'h58d : LOC <=          63'b000000000000000000000000000000000000000100000000000000100000000; // D (0x0000000000800100) 
    12'hace : LOC <=          63'b000000000000000000000000000000000000000100000000000001000000000; // D (0x0000000000800200) 
    12'h171 : LOC <=          63'b000000000000000000000000000000000000000100000000000010000000000; // D (0x0000000000800400) 
    12'h336 : LOC <=          63'b000000000000000000000000000000000000000100000000000100000000000; // D (0x0000000000800800) 
    12'h7b8 : LOC <=          63'b000000000000000000000000000000000000000100000000001000000000000; // D (0x0000000000801000) 
    12'hea4 : LOC <=          63'b000000000000000000000000000000000000000100000000010000000000000; // D (0x0000000000802000) 
    12'h9a5 : LOC <=          63'b000000000000000000000000000000000000000100000000100000000000000; // D (0x0000000000804000) 
    12'h7a7 : LOC <=          63'b000000000000000000000000000000000000000100000001000000000000000; // D (0x0000000000808000) 
    12'he9a : LOC <=          63'b000000000000000000000000000000000000000100000010000000000000000; // D (0x0000000000810000) 
    12'h9d9 : LOC <=          63'b000000000000000000000000000000000000000100000100000000000000000; // D (0x0000000000820000) 
    12'h75f : LOC <=          63'b000000000000000000000000000000000000000100001000000000000000000; // D (0x0000000000840000) 
    12'hf6a : LOC <=          63'b000000000000000000000000000000000000000100010000000000000000000; // D (0x0000000000880000) 
    12'ha39 : LOC <=          63'b000000000000000000000000000000000000000100100000000000000000000; // D (0x0000000000900000) 
    12'h09f : LOC <=          63'b000000000000000000000000000000000000000101000000000000000000000; // D (0x0000000000a00000) 
    12'h0ea : LOC <=          63'b000000000000000000000000000000000000000110000000000000000000000; // D (0x0000000000c00000) 
    12'hc5b : LOC <=          63'b000000000000000000000000000000000000000100000000000000000000000; // S (0x0000000000800000) 
//    12'h1d4 : LOC <=          63'b000000000000000000000000000000000000001100000000000000000000000; // D (0x0000000001800000) 
//    12'h27c : LOC <=          63'b000000000000000000000000000000000000010100000000000000000000000; // D (0x0000000002800000) 
//    12'h52c : LOC <=          63'b000000000000000000000000000000000000100100000000000000000000000; // D (0x0000000004800000) 
//    12'hb8c : LOC <=          63'b000000000000000000000000000000000001000100000000000000000000000; // D (0x0000000008800000) 
//    12'h3f5 : LOC <=          63'b000000000000000000000000000000000010000100000000000000000000000; // D (0x0000000010800000) 
//    12'h63e : LOC <=          63'b000000000000000000000000000000000100000100000000000000000000000; // D (0x0000000020800000) 
//    12'hda8 : LOC <=          63'b000000000000000000000000000000001000000100000000000000000000000; // D (0x0000000040800000) 
//    12'hfbd : LOC <=          63'b000000000000000000000000000000010000000100000000000000000000000; // D (0x0000000080800000) 
//    12'hb97 : LOC <=          63'b000000000000000000000000000000100000000100000000000000000000000; // D (0x0000000100800000) 
//    12'h3c3 : LOC <=          63'b000000000000000000000000000001000000000100000000000000000000000; // D (0x0000000200800000) 
//    12'h652 : LOC <=          63'b000000000000000000000000000010000000000100000000000000000000000; // D (0x0000000400800000) 
//    12'hd70 : LOC <=          63'b000000000000000000000000000100000000000100000000000000000000000; // D (0x0000000800800000) 
//    12'he0d : LOC <=          63'b000000000000000000000000001000000000000100000000000000000000000; // D (0x0000001000800000) 
//    12'h8f7 : LOC <=          63'b000000000000000000000000010000000000000100000000000000000000000; // D (0x0000002000800000) 
//    12'h503 : LOC <=          63'b000000000000000000000000100000000000000100000000000000000000000; // D (0x0000004000800000) 
//    12'hbd2 : LOC <=          63'b000000000000000000000001000000000000000100000000000000000000000; // D (0x0000008000800000) 
//    12'h349 : LOC <=          63'b000000000000000000000010000000000000000100000000000000000000000; // D (0x0000010000800000) 
//    12'h746 : LOC <=          63'b000000000000000000000100000000000000000100000000000000000000000; // D (0x0000020000800000) 
//    12'hf58 : LOC <=          63'b000000000000000000001000000000000000000100000000000000000000000; // D (0x0000040000800000) 
//    12'ha5d : LOC <=          63'b000000000000000000010000000000000000000100000000000000000000000; // D (0x0000080000800000) 
//    12'h057 : LOC <=          63'b000000000000000000100000000000000000000100000000000000000000000; // D (0x0000100000800000) 
//    12'h17a : LOC <=          63'b000000000000000001000000000000000000000100000000000000000000000; // D (0x0000200000800000) 
//    12'h320 : LOC <=          63'b000000000000000010000000000000000000000100000000000000000000000; // D (0x0000400000800000) 
//    12'h794 : LOC <=          63'b000000000000000100000000000000000000000100000000000000000000000; // D (0x0000800000800000) 
//    12'hefc : LOC <=          63'b000000000000001000000000000000000000000100000000000000000000000; // D (0x0001000000800000) 
//    12'h915 : LOC <=          63'b000000000000010000000000000000000000000100000000000000000000000; // D (0x0002000000800000) 
//    12'h6c7 : LOC <=          63'b000000000000100000000000000000000000000100000000000000000000000; // D (0x0004000000800000) 
//    12'hc5a : LOC <=          63'b000000000001000000000000000000000000000100000000000000000000000; // D (0x0008000000800000) 
//    12'hc59 : LOC <=          63'b000000000010000000000000000000000000000100000000000000000000000; // D (0x0010000000800000) 
//    12'hc5f : LOC <=          63'b000000000100000000000000000000000000000100000000000000000000000; // D (0x0020000000800000) 
//    12'hc53 : LOC <=          63'b000000001000000000000000000000000000000100000000000000000000000; // D (0x0040000000800000) 
//    12'hc4b : LOC <=          63'b000000010000000000000000000000000000000100000000000000000000000; // D (0x0080000000800000) 
//    12'hc7b : LOC <=          63'b000000100000000000000000000000000000000100000000000000000000000; // D (0x0100000000800000) 
//    12'hc1b : LOC <=          63'b000001000000000000000000000000000000000100000000000000000000000; // D (0x0200000000800000) 
//    12'hcdb : LOC <=          63'b000010000000000000000000000000000000000100000000000000000000000; // D (0x0400000000800000) 
//    12'hd5b : LOC <=          63'b000100000000000000000000000000000000000100000000000000000000000; // D (0x0800000000800000) 
//    12'he5b : LOC <=          63'b001000000000000000000000000000000000000100000000000000000000000; // D (0x1000000000800000) 
//    12'h85b : LOC <=          63'b010000000000000000000000000000000000000100000000000000000000000; // D (0x2000000000800000) 
//    12'h45b : LOC <=          63'b100000000000000000000000000000000000000100000000000000000000000; // D (0x4000000000800000) 
    12'h8b6 : LOC <=          63'b000000000000000000000000000000000000001000000000000000000000001; // D (0x0000000001000001) 
    12'h7fd : LOC <=          63'b000000000000000000000000000000000000001000000000000000000000010; // D (0x0000000001000002) 
    12'hc52 : LOC <=          63'b000000000000000000000000000000000000001000000000000000000000100; // D (0x0000000001000004) 
    12'he35 : LOC <=          63'b000000000000000000000000000000000000001000000000000000000001000; // D (0x0000000001000008) 
    12'hafb : LOC <=          63'b000000000000000000000000000000000000001000000000000000000010000; // D (0x0000000001000010) 
    12'h367 : LOC <=          63'b000000000000000000000000000000000000001000000000000000000100000; // D (0x0000000001000020) 
    12'h566 : LOC <=          63'b000000000000000000000000000000000000001000000000000000001000000; // D (0x0000000001000040) 
    12'h964 : LOC <=          63'b000000000000000000000000000000000000001000000000000000010000000; // D (0x0000000001000080) 
    12'h459 : LOC <=          63'b000000000000000000000000000000000000001000000000000000100000000; // D (0x0000000001000100) 
    12'hb1a : LOC <=          63'b000000000000000000000000000000000000001000000000000001000000000; // D (0x0000000001000200) 
    12'h0a5 : LOC <=          63'b000000000000000000000000000000000000001000000000000010000000000; // D (0x0000000001000400) 
    12'h2e2 : LOC <=          63'b000000000000000000000000000000000000001000000000000100000000000; // D (0x0000000001000800) 
    12'h66c : LOC <=          63'b000000000000000000000000000000000000001000000000001000000000000; // D (0x0000000001001000) 
    12'hf70 : LOC <=          63'b000000000000000000000000000000000000001000000000010000000000000; // D (0x0000000001002000) 
    12'h871 : LOC <=          63'b000000000000000000000000000000000000001000000000100000000000000; // D (0x0000000001004000) 
    12'h673 : LOC <=          63'b000000000000000000000000000000000000001000000001000000000000000; // D (0x0000000001008000) 
    12'hf4e : LOC <=          63'b000000000000000000000000000000000000001000000010000000000000000; // D (0x0000000001010000) 
    12'h80d : LOC <=          63'b000000000000000000000000000000000000001000000100000000000000000; // D (0x0000000001020000) 
    12'h68b : LOC <=          63'b000000000000000000000000000000000000001000001000000000000000000; // D (0x0000000001040000) 
    12'hebe : LOC <=          63'b000000000000000000000000000000000000001000010000000000000000000; // D (0x0000000001080000) 
    12'hbed : LOC <=          63'b000000000000000000000000000000000000001000100000000000000000000; // D (0x0000000001100000) 
    12'h14b : LOC <=          63'b000000000000000000000000000000000000001001000000000000000000000; // D (0x0000000001200000) 
    12'h13e : LOC <=          63'b000000000000000000000000000000000000001010000000000000000000000; // D (0x0000000001400000) 
    12'h1d4 : LOC <=          63'b000000000000000000000000000000000000001100000000000000000000000; // D (0x0000000001800000) 
    12'hd8f : LOC <=          63'b000000000000000000000000000000000000001000000000000000000000000; // S (0x0000000001000000) 
//    12'h3a8 : LOC <=          63'b000000000000000000000000000000000000011000000000000000000000000; // D (0x0000000003000000) 
//    12'h4f8 : LOC <=          63'b000000000000000000000000000000000000101000000000000000000000000; // D (0x0000000005000000) 
//    12'ha58 : LOC <=          63'b000000000000000000000000000000000001001000000000000000000000000; // D (0x0000000009000000) 
//    12'h221 : LOC <=          63'b000000000000000000000000000000000010001000000000000000000000000; // D (0x0000000011000000) 
//    12'h7ea : LOC <=          63'b000000000000000000000000000000000100001000000000000000000000000; // D (0x0000000021000000) 
//    12'hc7c : LOC <=          63'b000000000000000000000000000000001000001000000000000000000000000; // D (0x0000000041000000) 
//    12'he69 : LOC <=          63'b000000000000000000000000000000010000001000000000000000000000000; // D (0x0000000081000000) 
//    12'ha43 : LOC <=          63'b000000000000000000000000000000100000001000000000000000000000000; // D (0x0000000101000000) 
//    12'h217 : LOC <=          63'b000000000000000000000000000001000000001000000000000000000000000; // D (0x0000000201000000) 
//    12'h786 : LOC <=          63'b000000000000000000000000000010000000001000000000000000000000000; // D (0x0000000401000000) 
//    12'hca4 : LOC <=          63'b000000000000000000000000000100000000001000000000000000000000000; // D (0x0000000801000000) 
//    12'hfd9 : LOC <=          63'b000000000000000000000000001000000000001000000000000000000000000; // D (0x0000001001000000) 
//    12'h923 : LOC <=          63'b000000000000000000000000010000000000001000000000000000000000000; // D (0x0000002001000000) 
//    12'h4d7 : LOC <=          63'b000000000000000000000000100000000000001000000000000000000000000; // D (0x0000004001000000) 
//    12'ha06 : LOC <=          63'b000000000000000000000001000000000000001000000000000000000000000; // D (0x0000008001000000) 
//    12'h29d : LOC <=          63'b000000000000000000000010000000000000001000000000000000000000000; // D (0x0000010001000000) 
//    12'h692 : LOC <=          63'b000000000000000000000100000000000000001000000000000000000000000; // D (0x0000020001000000) 
//    12'he8c : LOC <=          63'b000000000000000000001000000000000000001000000000000000000000000; // D (0x0000040001000000) 
//    12'hb89 : LOC <=          63'b000000000000000000010000000000000000001000000000000000000000000; // D (0x0000080001000000) 
//    12'h183 : LOC <=          63'b000000000000000000100000000000000000001000000000000000000000000; // D (0x0000100001000000) 
//    12'h0ae : LOC <=          63'b000000000000000001000000000000000000001000000000000000000000000; // D (0x0000200001000000) 
//    12'h2f4 : LOC <=          63'b000000000000000010000000000000000000001000000000000000000000000; // D (0x0000400001000000) 
//    12'h640 : LOC <=          63'b000000000000000100000000000000000000001000000000000000000000000; // D (0x0000800001000000) 
//    12'hf28 : LOC <=          63'b000000000000001000000000000000000000001000000000000000000000000; // D (0x0001000001000000) 
//    12'h8c1 : LOC <=          63'b000000000000010000000000000000000000001000000000000000000000000; // D (0x0002000001000000) 
//    12'h713 : LOC <=          63'b000000000000100000000000000000000000001000000000000000000000000; // D (0x0004000001000000) 
//    12'hd8e : LOC <=          63'b000000000001000000000000000000000000001000000000000000000000000; // D (0x0008000001000000) 
//    12'hd8d : LOC <=          63'b000000000010000000000000000000000000001000000000000000000000000; // D (0x0010000001000000) 
//    12'hd8b : LOC <=          63'b000000000100000000000000000000000000001000000000000000000000000; // D (0x0020000001000000) 
//    12'hd87 : LOC <=          63'b000000001000000000000000000000000000001000000000000000000000000; // D (0x0040000001000000) 
//    12'hd9f : LOC <=          63'b000000010000000000000000000000000000001000000000000000000000000; // D (0x0080000001000000) 
//    12'hdaf : LOC <=          63'b000000100000000000000000000000000000001000000000000000000000000; // D (0x0100000001000000) 
//    12'hdcf : LOC <=          63'b000001000000000000000000000000000000001000000000000000000000000; // D (0x0200000001000000) 
//    12'hd0f : LOC <=          63'b000010000000000000000000000000000000001000000000000000000000000; // D (0x0400000001000000) 
//    12'hc8f : LOC <=          63'b000100000000000000000000000000000000001000000000000000000000000; // D (0x0800000001000000) 
//    12'hf8f : LOC <=          63'b001000000000000000000000000000000000001000000000000000000000000; // D (0x1000000001000000) 
//    12'h98f : LOC <=          63'b010000000000000000000000000000000000001000000000000000000000000; // D (0x2000000001000000) 
//    12'h58f : LOC <=          63'b100000000000000000000000000000000000001000000000000000000000000; // D (0x4000000001000000) 
    12'hb1e : LOC <=          63'b000000000000000000000000000000000000010000000000000000000000001; // D (0x0000000002000001) 
    12'h455 : LOC <=          63'b000000000000000000000000000000000000010000000000000000000000010; // D (0x0000000002000002) 
    12'hffa : LOC <=          63'b000000000000000000000000000000000000010000000000000000000000100; // D (0x0000000002000004) 
    12'hd9d : LOC <=          63'b000000000000000000000000000000000000010000000000000000000001000; // D (0x0000000002000008) 
    12'h953 : LOC <=          63'b000000000000000000000000000000000000010000000000000000000010000; // D (0x0000000002000010) 
    12'h0cf : LOC <=          63'b000000000000000000000000000000000000010000000000000000000100000; // D (0x0000000002000020) 
    12'h6ce : LOC <=          63'b000000000000000000000000000000000000010000000000000000001000000; // D (0x0000000002000040) 
    12'hacc : LOC <=          63'b000000000000000000000000000000000000010000000000000000010000000; // D (0x0000000002000080) 
    12'h7f1 : LOC <=          63'b000000000000000000000000000000000000010000000000000000100000000; // D (0x0000000002000100) 
    12'h8b2 : LOC <=          63'b000000000000000000000000000000000000010000000000000001000000000; // D (0x0000000002000200) 
    12'h30d : LOC <=          63'b000000000000000000000000000000000000010000000000000010000000000; // D (0x0000000002000400) 
    12'h14a : LOC <=          63'b000000000000000000000000000000000000010000000000000100000000000; // D (0x0000000002000800) 
    12'h5c4 : LOC <=          63'b000000000000000000000000000000000000010000000000001000000000000; // D (0x0000000002001000) 
    12'hcd8 : LOC <=          63'b000000000000000000000000000000000000010000000000010000000000000; // D (0x0000000002002000) 
    12'hbd9 : LOC <=          63'b000000000000000000000000000000000000010000000000100000000000000; // D (0x0000000002004000) 
    12'h5db : LOC <=          63'b000000000000000000000000000000000000010000000001000000000000000; // D (0x0000000002008000) 
    12'hce6 : LOC <=          63'b000000000000000000000000000000000000010000000010000000000000000; // D (0x0000000002010000) 
    12'hba5 : LOC <=          63'b000000000000000000000000000000000000010000000100000000000000000; // D (0x0000000002020000) 
    12'h523 : LOC <=          63'b000000000000000000000000000000000000010000001000000000000000000; // D (0x0000000002040000) 
    12'hd16 : LOC <=          63'b000000000000000000000000000000000000010000010000000000000000000; // D (0x0000000002080000) 
    12'h845 : LOC <=          63'b000000000000000000000000000000000000010000100000000000000000000; // D (0x0000000002100000) 
    12'h2e3 : LOC <=          63'b000000000000000000000000000000000000010001000000000000000000000; // D (0x0000000002200000) 
    12'h296 : LOC <=          63'b000000000000000000000000000000000000010010000000000000000000000; // D (0x0000000002400000) 
    12'h27c : LOC <=          63'b000000000000000000000000000000000000010100000000000000000000000; // D (0x0000000002800000) 
    12'h3a8 : LOC <=          63'b000000000000000000000000000000000000011000000000000000000000000; // D (0x0000000003000000) 
    12'he27 : LOC <=          63'b000000000000000000000000000000000000010000000000000000000000000; // S (0x0000000002000000) 
//    12'h750 : LOC <=          63'b000000000000000000000000000000000000110000000000000000000000000; // D (0x0000000006000000) 
//    12'h9f0 : LOC <=          63'b000000000000000000000000000000000001010000000000000000000000000; // D (0x000000000a000000) 
//    12'h189 : LOC <=          63'b000000000000000000000000000000000010010000000000000000000000000; // D (0x0000000012000000) 
//    12'h442 : LOC <=          63'b000000000000000000000000000000000100010000000000000000000000000; // D (0x0000000022000000) 
//    12'hfd4 : LOC <=          63'b000000000000000000000000000000001000010000000000000000000000000; // D (0x0000000042000000) 
//    12'hdc1 : LOC <=          63'b000000000000000000000000000000010000010000000000000000000000000; // D (0x0000000082000000) 
//    12'h9eb : LOC <=          63'b000000000000000000000000000000100000010000000000000000000000000; // D (0x0000000102000000) 
//    12'h1bf : LOC <=          63'b000000000000000000000000000001000000010000000000000000000000000; // D (0x0000000202000000) 
//    12'h42e : LOC <=          63'b000000000000000000000000000010000000010000000000000000000000000; // D (0x0000000402000000) 
//    12'hf0c : LOC <=          63'b000000000000000000000000000100000000010000000000000000000000000; // D (0x0000000802000000) 
//    12'hc71 : LOC <=          63'b000000000000000000000000001000000000010000000000000000000000000; // D (0x0000001002000000) 
//    12'ha8b : LOC <=          63'b000000000000000000000000010000000000010000000000000000000000000; // D (0x0000002002000000) 
//    12'h77f : LOC <=          63'b000000000000000000000000100000000000010000000000000000000000000; // D (0x0000004002000000) 
//    12'h9ae : LOC <=          63'b000000000000000000000001000000000000010000000000000000000000000; // D (0x0000008002000000) 
//    12'h135 : LOC <=          63'b000000000000000000000010000000000000010000000000000000000000000; // D (0x0000010002000000) 
//    12'h53a : LOC <=          63'b000000000000000000000100000000000000010000000000000000000000000; // D (0x0000020002000000) 
//    12'hd24 : LOC <=          63'b000000000000000000001000000000000000010000000000000000000000000; // D (0x0000040002000000) 
//    12'h821 : LOC <=          63'b000000000000000000010000000000000000010000000000000000000000000; // D (0x0000080002000000) 
//    12'h22b : LOC <=          63'b000000000000000000100000000000000000010000000000000000000000000; // D (0x0000100002000000) 
//    12'h306 : LOC <=          63'b000000000000000001000000000000000000010000000000000000000000000; // D (0x0000200002000000) 
//    12'h15c : LOC <=          63'b000000000000000010000000000000000000010000000000000000000000000; // D (0x0000400002000000) 
//    12'h5e8 : LOC <=          63'b000000000000000100000000000000000000010000000000000000000000000; // D (0x0000800002000000) 
//    12'hc80 : LOC <=          63'b000000000000001000000000000000000000010000000000000000000000000; // D (0x0001000002000000) 
//    12'hb69 : LOC <=          63'b000000000000010000000000000000000000010000000000000000000000000; // D (0x0002000002000000) 
//    12'h4bb : LOC <=          63'b000000000000100000000000000000000000010000000000000000000000000; // D (0x0004000002000000) 
//    12'he26 : LOC <=          63'b000000000001000000000000000000000000010000000000000000000000000; // D (0x0008000002000000) 
//    12'he25 : LOC <=          63'b000000000010000000000000000000000000010000000000000000000000000; // D (0x0010000002000000) 
//    12'he23 : LOC <=          63'b000000000100000000000000000000000000010000000000000000000000000; // D (0x0020000002000000) 
//    12'he2f : LOC <=          63'b000000001000000000000000000000000000010000000000000000000000000; // D (0x0040000002000000) 
//    12'he37 : LOC <=          63'b000000010000000000000000000000000000010000000000000000000000000; // D (0x0080000002000000) 
//    12'he07 : LOC <=          63'b000000100000000000000000000000000000010000000000000000000000000; // D (0x0100000002000000) 
//    12'he67 : LOC <=          63'b000001000000000000000000000000000000010000000000000000000000000; // D (0x0200000002000000) 
//    12'hea7 : LOC <=          63'b000010000000000000000000000000000000010000000000000000000000000; // D (0x0400000002000000) 
//    12'hf27 : LOC <=          63'b000100000000000000000000000000000000010000000000000000000000000; // D (0x0800000002000000) 
//    12'hc27 : LOC <=          63'b001000000000000000000000000000000000010000000000000000000000000; // D (0x1000000002000000) 
//    12'ha27 : LOC <=          63'b010000000000000000000000000000000000010000000000000000000000000; // D (0x2000000002000000) 
//    12'h627 : LOC <=          63'b100000000000000000000000000000000000010000000000000000000000000; // D (0x4000000002000000) 
    12'hc4e : LOC <=          63'b000000000000000000000000000000000000100000000000000000000000001; // D (0x0000000004000001) 
    12'h305 : LOC <=          63'b000000000000000000000000000000000000100000000000000000000000010; // D (0x0000000004000002) 
    12'h8aa : LOC <=          63'b000000000000000000000000000000000000100000000000000000000000100; // D (0x0000000004000004) 
    12'hacd : LOC <=          63'b000000000000000000000000000000000000100000000000000000000001000; // D (0x0000000004000008) 
    12'he03 : LOC <=          63'b000000000000000000000000000000000000100000000000000000000010000; // D (0x0000000004000010) 
    12'h79f : LOC <=          63'b000000000000000000000000000000000000100000000000000000000100000; // D (0x0000000004000020) 
    12'h19e : LOC <=          63'b000000000000000000000000000000000000100000000000000000001000000; // D (0x0000000004000040) 
    12'hd9c : LOC <=          63'b000000000000000000000000000000000000100000000000000000010000000; // D (0x0000000004000080) 
    12'h0a1 : LOC <=          63'b000000000000000000000000000000000000100000000000000000100000000; // D (0x0000000004000100) 
    12'hfe2 : LOC <=          63'b000000000000000000000000000000000000100000000000000001000000000; // D (0x0000000004000200) 
    12'h45d : LOC <=          63'b000000000000000000000000000000000000100000000000000010000000000; // D (0x0000000004000400) 
    12'h61a : LOC <=          63'b000000000000000000000000000000000000100000000000000100000000000; // D (0x0000000004000800) 
    12'h294 : LOC <=          63'b000000000000000000000000000000000000100000000000001000000000000; // D (0x0000000004001000) 
    12'hb88 : LOC <=          63'b000000000000000000000000000000000000100000000000010000000000000; // D (0x0000000004002000) 
    12'hc89 : LOC <=          63'b000000000000000000000000000000000000100000000000100000000000000; // D (0x0000000004004000) 
    12'h28b : LOC <=          63'b000000000000000000000000000000000000100000000001000000000000000; // D (0x0000000004008000) 
    12'hbb6 : LOC <=          63'b000000000000000000000000000000000000100000000010000000000000000; // D (0x0000000004010000) 
    12'hcf5 : LOC <=          63'b000000000000000000000000000000000000100000000100000000000000000; // D (0x0000000004020000) 
    12'h273 : LOC <=          63'b000000000000000000000000000000000000100000001000000000000000000; // D (0x0000000004040000) 
    12'ha46 : LOC <=          63'b000000000000000000000000000000000000100000010000000000000000000; // D (0x0000000004080000) 
    12'hf15 : LOC <=          63'b000000000000000000000000000000000000100000100000000000000000000; // D (0x0000000004100000) 
    12'h5b3 : LOC <=          63'b000000000000000000000000000000000000100001000000000000000000000; // D (0x0000000004200000) 
    12'h5c6 : LOC <=          63'b000000000000000000000000000000000000100010000000000000000000000; // D (0x0000000004400000) 
    12'h52c : LOC <=          63'b000000000000000000000000000000000000100100000000000000000000000; // D (0x0000000004800000) 
    12'h4f8 : LOC <=          63'b000000000000000000000000000000000000101000000000000000000000000; // D (0x0000000005000000) 
    12'h750 : LOC <=          63'b000000000000000000000000000000000000110000000000000000000000000; // D (0x0000000006000000) 
    12'h977 : LOC <=          63'b000000000000000000000000000000000000100000000000000000000000000; // S (0x0000000004000000) 
//    12'hea0 : LOC <=          63'b000000000000000000000000000000000001100000000000000000000000000; // D (0x000000000c000000) 
//    12'h6d9 : LOC <=          63'b000000000000000000000000000000000010100000000000000000000000000; // D (0x0000000014000000) 
//    12'h312 : LOC <=          63'b000000000000000000000000000000000100100000000000000000000000000; // D (0x0000000024000000) 
//    12'h884 : LOC <=          63'b000000000000000000000000000000001000100000000000000000000000000; // D (0x0000000044000000) 
//    12'ha91 : LOC <=          63'b000000000000000000000000000000010000100000000000000000000000000; // D (0x0000000084000000) 
//    12'hebb : LOC <=          63'b000000000000000000000000000000100000100000000000000000000000000; // D (0x0000000104000000) 
//    12'h6ef : LOC <=          63'b000000000000000000000000000001000000100000000000000000000000000; // D (0x0000000204000000) 
//    12'h37e : LOC <=          63'b000000000000000000000000000010000000100000000000000000000000000; // D (0x0000000404000000) 
//    12'h85c : LOC <=          63'b000000000000000000000000000100000000100000000000000000000000000; // D (0x0000000804000000) 
//    12'hb21 : LOC <=          63'b000000000000000000000000001000000000100000000000000000000000000; // D (0x0000001004000000) 
//    12'hddb : LOC <=          63'b000000000000000000000000010000000000100000000000000000000000000; // D (0x0000002004000000) 
//    12'h02f : LOC <=          63'b000000000000000000000000100000000000100000000000000000000000000; // D (0x0000004004000000) 
//    12'hefe : LOC <=          63'b000000000000000000000001000000000000100000000000000000000000000; // D (0x0000008004000000) 
//    12'h665 : LOC <=          63'b000000000000000000000010000000000000100000000000000000000000000; // D (0x0000010004000000) 
//    12'h26a : LOC <=          63'b000000000000000000000100000000000000100000000000000000000000000; // D (0x0000020004000000) 
//    12'ha74 : LOC <=          63'b000000000000000000001000000000000000100000000000000000000000000; // D (0x0000040004000000) 
//    12'hf71 : LOC <=          63'b000000000000000000010000000000000000100000000000000000000000000; // D (0x0000080004000000) 
//    12'h57b : LOC <=          63'b000000000000000000100000000000000000100000000000000000000000000; // D (0x0000100004000000) 
//    12'h456 : LOC <=          63'b000000000000000001000000000000000000100000000000000000000000000; // D (0x0000200004000000) 
//    12'h60c : LOC <=          63'b000000000000000010000000000000000000100000000000000000000000000; // D (0x0000400004000000) 
//    12'h2b8 : LOC <=          63'b000000000000000100000000000000000000100000000000000000000000000; // D (0x0000800004000000) 
//    12'hbd0 : LOC <=          63'b000000000000001000000000000000000000100000000000000000000000000; // D (0x0001000004000000) 
//    12'hc39 : LOC <=          63'b000000000000010000000000000000000000100000000000000000000000000; // D (0x0002000004000000) 
//    12'h3eb : LOC <=          63'b000000000000100000000000000000000000100000000000000000000000000; // D (0x0004000004000000) 
//    12'h976 : LOC <=          63'b000000000001000000000000000000000000100000000000000000000000000; // D (0x0008000004000000) 
//    12'h975 : LOC <=          63'b000000000010000000000000000000000000100000000000000000000000000; // D (0x0010000004000000) 
//    12'h973 : LOC <=          63'b000000000100000000000000000000000000100000000000000000000000000; // D (0x0020000004000000) 
//    12'h97f : LOC <=          63'b000000001000000000000000000000000000100000000000000000000000000; // D (0x0040000004000000) 
//    12'h967 : LOC <=          63'b000000010000000000000000000000000000100000000000000000000000000; // D (0x0080000004000000) 
//    12'h957 : LOC <=          63'b000000100000000000000000000000000000100000000000000000000000000; // D (0x0100000004000000) 
//    12'h937 : LOC <=          63'b000001000000000000000000000000000000100000000000000000000000000; // D (0x0200000004000000) 
//    12'h9f7 : LOC <=          63'b000010000000000000000000000000000000100000000000000000000000000; // D (0x0400000004000000) 
//    12'h877 : LOC <=          63'b000100000000000000000000000000000000100000000000000000000000000; // D (0x0800000004000000) 
//    12'hb77 : LOC <=          63'b001000000000000000000000000000000000100000000000000000000000000; // D (0x1000000004000000) 
//    12'hd77 : LOC <=          63'b010000000000000000000000000000000000100000000000000000000000000; // D (0x2000000004000000) 
//    12'h177 : LOC <=          63'b100000000000000000000000000000000000100000000000000000000000000; // D (0x4000000004000000) 
    12'h2ee : LOC <=          63'b000000000000000000000000000000000001000000000000000000000000001; // D (0x0000000008000001) 
    12'hda5 : LOC <=          63'b000000000000000000000000000000000001000000000000000000000000010; // D (0x0000000008000002) 
    12'h60a : LOC <=          63'b000000000000000000000000000000000001000000000000000000000000100; // D (0x0000000008000004) 
    12'h46d : LOC <=          63'b000000000000000000000000000000000001000000000000000000000001000; // D (0x0000000008000008) 
    12'h0a3 : LOC <=          63'b000000000000000000000000000000000001000000000000000000000010000; // D (0x0000000008000010) 
    12'h93f : LOC <=          63'b000000000000000000000000000000000001000000000000000000000100000; // D (0x0000000008000020) 
    12'hf3e : LOC <=          63'b000000000000000000000000000000000001000000000000000000001000000; // D (0x0000000008000040) 
    12'h33c : LOC <=          63'b000000000000000000000000000000000001000000000000000000010000000; // D (0x0000000008000080) 
    12'he01 : LOC <=          63'b000000000000000000000000000000000001000000000000000000100000000; // D (0x0000000008000100) 
    12'h142 : LOC <=          63'b000000000000000000000000000000000001000000000000000001000000000; // D (0x0000000008000200) 
    12'hafd : LOC <=          63'b000000000000000000000000000000000001000000000000000010000000000; // D (0x0000000008000400) 
    12'h8ba : LOC <=          63'b000000000000000000000000000000000001000000000000000100000000000; // D (0x0000000008000800) 
    12'hc34 : LOC <=          63'b000000000000000000000000000000000001000000000000001000000000000; // D (0x0000000008001000) 
    12'h528 : LOC <=          63'b000000000000000000000000000000000001000000000000010000000000000; // D (0x0000000008002000) 
    12'h229 : LOC <=          63'b000000000000000000000000000000000001000000000000100000000000000; // D (0x0000000008004000) 
    12'hc2b : LOC <=          63'b000000000000000000000000000000000001000000000001000000000000000; // D (0x0000000008008000) 
    12'h516 : LOC <=          63'b000000000000000000000000000000000001000000000010000000000000000; // D (0x0000000008010000) 
    12'h255 : LOC <=          63'b000000000000000000000000000000000001000000000100000000000000000; // D (0x0000000008020000) 
    12'hcd3 : LOC <=          63'b000000000000000000000000000000000001000000001000000000000000000; // D (0x0000000008040000) 
    12'h4e6 : LOC <=          63'b000000000000000000000000000000000001000000010000000000000000000; // D (0x0000000008080000) 
    12'h1b5 : LOC <=          63'b000000000000000000000000000000000001000000100000000000000000000; // D (0x0000000008100000) 
    12'hb13 : LOC <=          63'b000000000000000000000000000000000001000001000000000000000000000; // D (0x0000000008200000) 
    12'hb66 : LOC <=          63'b000000000000000000000000000000000001000010000000000000000000000; // D (0x0000000008400000) 
    12'hb8c : LOC <=          63'b000000000000000000000000000000000001000100000000000000000000000; // D (0x0000000008800000) 
    12'ha58 : LOC <=          63'b000000000000000000000000000000000001001000000000000000000000000; // D (0x0000000009000000) 
    12'h9f0 : LOC <=          63'b000000000000000000000000000000000001010000000000000000000000000; // D (0x000000000a000000) 
    12'hea0 : LOC <=          63'b000000000000000000000000000000000001100000000000000000000000000; // D (0x000000000c000000) 
    12'h7d7 : LOC <=          63'b000000000000000000000000000000000001000000000000000000000000000; // S (0x0000000008000000) 
//    12'h879 : LOC <=          63'b000000000000000000000000000000000011000000000000000000000000000; // D (0x0000000018000000) 
//    12'hdb2 : LOC <=          63'b000000000000000000000000000000000101000000000000000000000000000; // D (0x0000000028000000) 
//    12'h624 : LOC <=          63'b000000000000000000000000000000001001000000000000000000000000000; // D (0x0000000048000000) 
//    12'h431 : LOC <=          63'b000000000000000000000000000000010001000000000000000000000000000; // D (0x0000000088000000) 
//    12'h01b : LOC <=          63'b000000000000000000000000000000100001000000000000000000000000000; // D (0x0000000108000000) 
//    12'h84f : LOC <=          63'b000000000000000000000000000001000001000000000000000000000000000; // D (0x0000000208000000) 
//    12'hdde : LOC <=          63'b000000000000000000000000000010000001000000000000000000000000000; // D (0x0000000408000000) 
//    12'h6fc : LOC <=          63'b000000000000000000000000000100000001000000000000000000000000000; // D (0x0000000808000000) 
//    12'h581 : LOC <=          63'b000000000000000000000000001000000001000000000000000000000000000; // D (0x0000001008000000) 
//    12'h37b : LOC <=          63'b000000000000000000000000010000000001000000000000000000000000000; // D (0x0000002008000000) 
//    12'he8f : LOC <=          63'b000000000000000000000000100000000001000000000000000000000000000; // D (0x0000004008000000) 
//    12'h05e : LOC <=          63'b000000000000000000000001000000000001000000000000000000000000000; // D (0x0000008008000000) 
//    12'h8c5 : LOC <=          63'b000000000000000000000010000000000001000000000000000000000000000; // D (0x0000010008000000) 
//    12'hcca : LOC <=          63'b000000000000000000000100000000000001000000000000000000000000000; // D (0x0000020008000000) 
//    12'h4d4 : LOC <=          63'b000000000000000000001000000000000001000000000000000000000000000; // D (0x0000040008000000) 
//    12'h1d1 : LOC <=          63'b000000000000000000010000000000000001000000000000000000000000000; // D (0x0000080008000000) 
//    12'hbdb : LOC <=          63'b000000000000000000100000000000000001000000000000000000000000000; // D (0x0000100008000000) 
//    12'haf6 : LOC <=          63'b000000000000000001000000000000000001000000000000000000000000000; // D (0x0000200008000000) 
//    12'h8ac : LOC <=          63'b000000000000000010000000000000000001000000000000000000000000000; // D (0x0000400008000000) 
//    12'hc18 : LOC <=          63'b000000000000000100000000000000000001000000000000000000000000000; // D (0x0000800008000000) 
//    12'h570 : LOC <=          63'b000000000000001000000000000000000001000000000000000000000000000; // D (0x0001000008000000) 
//    12'h299 : LOC <=          63'b000000000000010000000000000000000001000000000000000000000000000; // D (0x0002000008000000) 
//    12'hd4b : LOC <=          63'b000000000000100000000000000000000001000000000000000000000000000; // D (0x0004000008000000) 
//    12'h7d6 : LOC <=          63'b000000000001000000000000000000000001000000000000000000000000000; // D (0x0008000008000000) 
//    12'h7d5 : LOC <=          63'b000000000010000000000000000000000001000000000000000000000000000; // D (0x0010000008000000) 
//    12'h7d3 : LOC <=          63'b000000000100000000000000000000000001000000000000000000000000000; // D (0x0020000008000000) 
//    12'h7df : LOC <=          63'b000000001000000000000000000000000001000000000000000000000000000; // D (0x0040000008000000) 
//    12'h7c7 : LOC <=          63'b000000010000000000000000000000000001000000000000000000000000000; // D (0x0080000008000000) 
//    12'h7f7 : LOC <=          63'b000000100000000000000000000000000001000000000000000000000000000; // D (0x0100000008000000) 
//    12'h797 : LOC <=          63'b000001000000000000000000000000000001000000000000000000000000000; // D (0x0200000008000000) 
//    12'h757 : LOC <=          63'b000010000000000000000000000000000001000000000000000000000000000; // D (0x0400000008000000) 
//    12'h6d7 : LOC <=          63'b000100000000000000000000000000000001000000000000000000000000000; // D (0x0800000008000000) 
//    12'h5d7 : LOC <=          63'b001000000000000000000000000000000001000000000000000000000000000; // D (0x1000000008000000) 
//    12'h3d7 : LOC <=          63'b010000000000000000000000000000000001000000000000000000000000000; // D (0x2000000008000000) 
//    12'hfd7 : LOC <=          63'b100000000000000000000000000000000001000000000000000000000000000; // D (0x4000000008000000) 
    12'ha97 : LOC <=          63'b000000000000000000000000000000000010000000000000000000000000001; // D (0x0000000010000001) 
    12'h5dc : LOC <=          63'b000000000000000000000000000000000010000000000000000000000000010; // D (0x0000000010000002) 
    12'he73 : LOC <=          63'b000000000000000000000000000000000010000000000000000000000000100; // D (0x0000000010000004) 
    12'hc14 : LOC <=          63'b000000000000000000000000000000000010000000000000000000000001000; // D (0x0000000010000008) 
    12'h8da : LOC <=          63'b000000000000000000000000000000000010000000000000000000000010000; // D (0x0000000010000010) 
    12'h146 : LOC <=          63'b000000000000000000000000000000000010000000000000000000000100000; // D (0x0000000010000020) 
    12'h747 : LOC <=          63'b000000000000000000000000000000000010000000000000000000001000000; // D (0x0000000010000040) 
    12'hb45 : LOC <=          63'b000000000000000000000000000000000010000000000000000000010000000; // D (0x0000000010000080) 
    12'h678 : LOC <=          63'b000000000000000000000000000000000010000000000000000000100000000; // D (0x0000000010000100) 
    12'h93b : LOC <=          63'b000000000000000000000000000000000010000000000000000001000000000; // D (0x0000000010000200) 
    12'h284 : LOC <=          63'b000000000000000000000000000000000010000000000000000010000000000; // D (0x0000000010000400) 
    12'h0c3 : LOC <=          63'b000000000000000000000000000000000010000000000000000100000000000; // D (0x0000000010000800) 
    12'h44d : LOC <=          63'b000000000000000000000000000000000010000000000000001000000000000; // D (0x0000000010001000) 
    12'hd51 : LOC <=          63'b000000000000000000000000000000000010000000000000010000000000000; // D (0x0000000010002000) 
    12'ha50 : LOC <=          63'b000000000000000000000000000000000010000000000000100000000000000; // D (0x0000000010004000) 
    12'h452 : LOC <=          63'b000000000000000000000000000000000010000000000001000000000000000; // D (0x0000000010008000) 
    12'hd6f : LOC <=          63'b000000000000000000000000000000000010000000000010000000000000000; // D (0x0000000010010000) 
    12'ha2c : LOC <=          63'b000000000000000000000000000000000010000000000100000000000000000; // D (0x0000000010020000) 
    12'h4aa : LOC <=          63'b000000000000000000000000000000000010000000001000000000000000000; // D (0x0000000010040000) 
    12'hc9f : LOC <=          63'b000000000000000000000000000000000010000000010000000000000000000; // D (0x0000000010080000) 
    12'h9cc : LOC <=          63'b000000000000000000000000000000000010000000100000000000000000000; // D (0x0000000010100000) 
    12'h36a : LOC <=          63'b000000000000000000000000000000000010000001000000000000000000000; // D (0x0000000010200000) 
    12'h31f : LOC <=          63'b000000000000000000000000000000000010000010000000000000000000000; // D (0x0000000010400000) 
    12'h3f5 : LOC <=          63'b000000000000000000000000000000000010000100000000000000000000000; // D (0x0000000010800000) 
    12'h221 : LOC <=          63'b000000000000000000000000000000000010001000000000000000000000000; // D (0x0000000011000000) 
    12'h189 : LOC <=          63'b000000000000000000000000000000000010010000000000000000000000000; // D (0x0000000012000000) 
    12'h6d9 : LOC <=          63'b000000000000000000000000000000000010100000000000000000000000000; // D (0x0000000014000000) 
    12'h879 : LOC <=          63'b000000000000000000000000000000000011000000000000000000000000000; // D (0x0000000018000000) 
    12'hfae : LOC <=          63'b000000000000000000000000000000000010000000000000000000000000000; // S (0x0000000010000000) 
//    12'h5cb : LOC <=          63'b000000000000000000000000000000000110000000000000000000000000000; // D (0x0000000030000000) 
//    12'he5d : LOC <=          63'b000000000000000000000000000000001010000000000000000000000000000; // D (0x0000000050000000) 
//    12'hc48 : LOC <=          63'b000000000000000000000000000000010010000000000000000000000000000; // D (0x0000000090000000) 
//    12'h862 : LOC <=          63'b000000000000000000000000000000100010000000000000000000000000000; // D (0x0000000110000000) 
//    12'h036 : LOC <=          63'b000000000000000000000000000001000010000000000000000000000000000; // D (0x0000000210000000) 
//    12'h5a7 : LOC <=          63'b000000000000000000000000000010000010000000000000000000000000000; // D (0x0000000410000000) 
//    12'he85 : LOC <=          63'b000000000000000000000000000100000010000000000000000000000000000; // D (0x0000000810000000) 
//    12'hdf8 : LOC <=          63'b000000000000000000000000001000000010000000000000000000000000000; // D (0x0000001010000000) 
//    12'hb02 : LOC <=          63'b000000000000000000000000010000000010000000000000000000000000000; // D (0x0000002010000000) 
//    12'h6f6 : LOC <=          63'b000000000000000000000000100000000010000000000000000000000000000; // D (0x0000004010000000) 
//    12'h827 : LOC <=          63'b000000000000000000000001000000000010000000000000000000000000000; // D (0x0000008010000000) 
//    12'h0bc : LOC <=          63'b000000000000000000000010000000000010000000000000000000000000000; // D (0x0000010010000000) 
//    12'h4b3 : LOC <=          63'b000000000000000000000100000000000010000000000000000000000000000; // D (0x0000020010000000) 
//    12'hcad : LOC <=          63'b000000000000000000001000000000000010000000000000000000000000000; // D (0x0000040010000000) 
//    12'h9a8 : LOC <=          63'b000000000000000000010000000000000010000000000000000000000000000; // D (0x0000080010000000) 
//    12'h3a2 : LOC <=          63'b000000000000000000100000000000000010000000000000000000000000000; // D (0x0000100010000000) 
//    12'h28f : LOC <=          63'b000000000000000001000000000000000010000000000000000000000000000; // D (0x0000200010000000) 
//    12'h0d5 : LOC <=          63'b000000000000000010000000000000000010000000000000000000000000000; // D (0x0000400010000000) 
//    12'h461 : LOC <=          63'b000000000000000100000000000000000010000000000000000000000000000; // D (0x0000800010000000) 
//    12'hd09 : LOC <=          63'b000000000000001000000000000000000010000000000000000000000000000; // D (0x0001000010000000) 
//    12'hae0 : LOC <=          63'b000000000000010000000000000000000010000000000000000000000000000; // D (0x0002000010000000) 
//    12'h532 : LOC <=          63'b000000000000100000000000000000000010000000000000000000000000000; // D (0x0004000010000000) 
//    12'hfaf : LOC <=          63'b000000000001000000000000000000000010000000000000000000000000000; // D (0x0008000010000000) 
//    12'hfac : LOC <=          63'b000000000010000000000000000000000010000000000000000000000000000; // D (0x0010000010000000) 
//    12'hfaa : LOC <=          63'b000000000100000000000000000000000010000000000000000000000000000; // D (0x0020000010000000) 
//    12'hfa6 : LOC <=          63'b000000001000000000000000000000000010000000000000000000000000000; // D (0x0040000010000000) 
//    12'hfbe : LOC <=          63'b000000010000000000000000000000000010000000000000000000000000000; // D (0x0080000010000000) 
//    12'hf8e : LOC <=          63'b000000100000000000000000000000000010000000000000000000000000000; // D (0x0100000010000000) 
//    12'hfee : LOC <=          63'b000001000000000000000000000000000010000000000000000000000000000; // D (0x0200000010000000) 
//    12'hf2e : LOC <=          63'b000010000000000000000000000000000010000000000000000000000000000; // D (0x0400000010000000) 
//    12'heae : LOC <=          63'b000100000000000000000000000000000010000000000000000000000000000; // D (0x0800000010000000) 
//    12'hdae : LOC <=          63'b001000000000000000000000000000000010000000000000000000000000000; // D (0x1000000010000000) 
//    12'hbae : LOC <=          63'b010000000000000000000000000000000010000000000000000000000000000; // D (0x2000000010000000) 
//    12'h7ae : LOC <=          63'b100000000000000000000000000000000010000000000000000000000000000; // D (0x4000000010000000) 
    12'hf5c : LOC <=          63'b000000000000000000000000000000000100000000000000000000000000001; // D (0x0000000020000001) 
    12'h017 : LOC <=          63'b000000000000000000000000000000000100000000000000000000000000010; // D (0x0000000020000002) 
    12'hbb8 : LOC <=          63'b000000000000000000000000000000000100000000000000000000000000100; // D (0x0000000020000004) 
    12'h9df : LOC <=          63'b000000000000000000000000000000000100000000000000000000000001000; // D (0x0000000020000008) 
    12'hd11 : LOC <=          63'b000000000000000000000000000000000100000000000000000000000010000; // D (0x0000000020000010) 
    12'h48d : LOC <=          63'b000000000000000000000000000000000100000000000000000000000100000; // D (0x0000000020000020) 
    12'h28c : LOC <=          63'b000000000000000000000000000000000100000000000000000000001000000; // D (0x0000000020000040) 
    12'he8e : LOC <=          63'b000000000000000000000000000000000100000000000000000000010000000; // D (0x0000000020000080) 
    12'h3b3 : LOC <=          63'b000000000000000000000000000000000100000000000000000000100000000; // D (0x0000000020000100) 
    12'hcf0 : LOC <=          63'b000000000000000000000000000000000100000000000000000001000000000; // D (0x0000000020000200) 
    12'h74f : LOC <=          63'b000000000000000000000000000000000100000000000000000010000000000; // D (0x0000000020000400) 
    12'h508 : LOC <=          63'b000000000000000000000000000000000100000000000000000100000000000; // D (0x0000000020000800) 
    12'h186 : LOC <=          63'b000000000000000000000000000000000100000000000000001000000000000; // D (0x0000000020001000) 
    12'h89a : LOC <=          63'b000000000000000000000000000000000100000000000000010000000000000; // D (0x0000000020002000) 
    12'hf9b : LOC <=          63'b000000000000000000000000000000000100000000000000100000000000000; // D (0x0000000020004000) 
    12'h199 : LOC <=          63'b000000000000000000000000000000000100000000000001000000000000000; // D (0x0000000020008000) 
    12'h8a4 : LOC <=          63'b000000000000000000000000000000000100000000000010000000000000000; // D (0x0000000020010000) 
    12'hfe7 : LOC <=          63'b000000000000000000000000000000000100000000000100000000000000000; // D (0x0000000020020000) 
    12'h161 : LOC <=          63'b000000000000000000000000000000000100000000001000000000000000000; // D (0x0000000020040000) 
    12'h954 : LOC <=          63'b000000000000000000000000000000000100000000010000000000000000000; // D (0x0000000020080000) 
    12'hc07 : LOC <=          63'b000000000000000000000000000000000100000000100000000000000000000; // D (0x0000000020100000) 
    12'h6a1 : LOC <=          63'b000000000000000000000000000000000100000001000000000000000000000; // D (0x0000000020200000) 
    12'h6d4 : LOC <=          63'b000000000000000000000000000000000100000010000000000000000000000; // D (0x0000000020400000) 
    12'h63e : LOC <=          63'b000000000000000000000000000000000100000100000000000000000000000; // D (0x0000000020800000) 
    12'h7ea : LOC <=          63'b000000000000000000000000000000000100001000000000000000000000000; // D (0x0000000021000000) 
    12'h442 : LOC <=          63'b000000000000000000000000000000000100010000000000000000000000000; // D (0x0000000022000000) 
    12'h312 : LOC <=          63'b000000000000000000000000000000000100100000000000000000000000000; // D (0x0000000024000000) 
    12'hdb2 : LOC <=          63'b000000000000000000000000000000000101000000000000000000000000000; // D (0x0000000028000000) 
    12'h5cb : LOC <=          63'b000000000000000000000000000000000110000000000000000000000000000; // D (0x0000000030000000) 
    12'ha65 : LOC <=          63'b000000000000000000000000000000000100000000000000000000000000000; // S (0x0000000020000000) 
//    12'hb96 : LOC <=          63'b000000000000000000000000000000001100000000000000000000000000000; // D (0x0000000060000000) 
//    12'h983 : LOC <=          63'b000000000000000000000000000000010100000000000000000000000000000; // D (0x00000000a0000000) 
//    12'hda9 : LOC <=          63'b000000000000000000000000000000100100000000000000000000000000000; // D (0x0000000120000000) 
//    12'h5fd : LOC <=          63'b000000000000000000000000000001000100000000000000000000000000000; // D (0x0000000220000000) 
//    12'h06c : LOC <=          63'b000000000000000000000000000010000100000000000000000000000000000; // D (0x0000000420000000) 
//    12'hb4e : LOC <=          63'b000000000000000000000000000100000100000000000000000000000000000; // D (0x0000000820000000) 
//    12'h833 : LOC <=          63'b000000000000000000000000001000000100000000000000000000000000000; // D (0x0000001020000000) 
//    12'hec9 : LOC <=          63'b000000000000000000000000010000000100000000000000000000000000000; // D (0x0000002020000000) 
//    12'h33d : LOC <=          63'b000000000000000000000000100000000100000000000000000000000000000; // D (0x0000004020000000) 
//    12'hdec : LOC <=          63'b000000000000000000000001000000000100000000000000000000000000000; // D (0x0000008020000000) 
//    12'h577 : LOC <=          63'b000000000000000000000010000000000100000000000000000000000000000; // D (0x0000010020000000) 
//    12'h178 : LOC <=          63'b000000000000000000000100000000000100000000000000000000000000000; // D (0x0000020020000000) 
//    12'h966 : LOC <=          63'b000000000000000000001000000000000100000000000000000000000000000; // D (0x0000040020000000) 
//    12'hc63 : LOC <=          63'b000000000000000000010000000000000100000000000000000000000000000; // D (0x0000080020000000) 
//    12'h669 : LOC <=          63'b000000000000000000100000000000000100000000000000000000000000000; // D (0x0000100020000000) 
//    12'h744 : LOC <=          63'b000000000000000001000000000000000100000000000000000000000000000; // D (0x0000200020000000) 
//    12'h51e : LOC <=          63'b000000000000000010000000000000000100000000000000000000000000000; // D (0x0000400020000000) 
//    12'h1aa : LOC <=          63'b000000000000000100000000000000000100000000000000000000000000000; // D (0x0000800020000000) 
//    12'h8c2 : LOC <=          63'b000000000000001000000000000000000100000000000000000000000000000; // D (0x0001000020000000) 
//    12'hf2b : LOC <=          63'b000000000000010000000000000000000100000000000000000000000000000; // D (0x0002000020000000) 
//    12'h0f9 : LOC <=          63'b000000000000100000000000000000000100000000000000000000000000000; // D (0x0004000020000000) 
//    12'ha64 : LOC <=          63'b000000000001000000000000000000000100000000000000000000000000000; // D (0x0008000020000000) 
//    12'ha67 : LOC <=          63'b000000000010000000000000000000000100000000000000000000000000000; // D (0x0010000020000000) 
//    12'ha61 : LOC <=          63'b000000000100000000000000000000000100000000000000000000000000000; // D (0x0020000020000000) 
//    12'ha6d : LOC <=          63'b000000001000000000000000000000000100000000000000000000000000000; // D (0x0040000020000000) 
//    12'ha75 : LOC <=          63'b000000010000000000000000000000000100000000000000000000000000000; // D (0x0080000020000000) 
//    12'ha45 : LOC <=          63'b000000100000000000000000000000000100000000000000000000000000000; // D (0x0100000020000000) 
//    12'ha25 : LOC <=          63'b000001000000000000000000000000000100000000000000000000000000000; // D (0x0200000020000000) 
//    12'hae5 : LOC <=          63'b000010000000000000000000000000000100000000000000000000000000000; // D (0x0400000020000000) 
//    12'hb65 : LOC <=          63'b000100000000000000000000000000000100000000000000000000000000000; // D (0x0800000020000000) 
//    12'h865 : LOC <=          63'b001000000000000000000000000000000100000000000000000000000000000; // D (0x1000000020000000) 
//    12'he65 : LOC <=          63'b010000000000000000000000000000000100000000000000000000000000000; // D (0x2000000020000000) 
//    12'h265 : LOC <=          63'b100000000000000000000000000000000100000000000000000000000000000; // D (0x4000000020000000) 
    12'h4ca : LOC <=          63'b000000000000000000000000000000001000000000000000000000000000001; // D (0x0000000040000001) 
    12'hb81 : LOC <=          63'b000000000000000000000000000000001000000000000000000000000000010; // D (0x0000000040000002) 
    12'h02e : LOC <=          63'b000000000000000000000000000000001000000000000000000000000000100; // D (0x0000000040000004) 
    12'h249 : LOC <=          63'b000000000000000000000000000000001000000000000000000000000001000; // D (0x0000000040000008) 
    12'h687 : LOC <=          63'b000000000000000000000000000000001000000000000000000000000010000; // D (0x0000000040000010) 
    12'hf1b : LOC <=          63'b000000000000000000000000000000001000000000000000000000000100000; // D (0x0000000040000020) 
    12'h91a : LOC <=          63'b000000000000000000000000000000001000000000000000000000001000000; // D (0x0000000040000040) 
    12'h518 : LOC <=          63'b000000000000000000000000000000001000000000000000000000010000000; // D (0x0000000040000080) 
    12'h825 : LOC <=          63'b000000000000000000000000000000001000000000000000000000100000000; // D (0x0000000040000100) 
    12'h766 : LOC <=          63'b000000000000000000000000000000001000000000000000000001000000000; // D (0x0000000040000200) 
    12'hcd9 : LOC <=          63'b000000000000000000000000000000001000000000000000000010000000000; // D (0x0000000040000400) 
    12'he9e : LOC <=          63'b000000000000000000000000000000001000000000000000000100000000000; // D (0x0000000040000800) 
    12'ha10 : LOC <=          63'b000000000000000000000000000000001000000000000000001000000000000; // D (0x0000000040001000) 
    12'h30c : LOC <=          63'b000000000000000000000000000000001000000000000000010000000000000; // D (0x0000000040002000) 
    12'h40d : LOC <=          63'b000000000000000000000000000000001000000000000000100000000000000; // D (0x0000000040004000) 
    12'ha0f : LOC <=          63'b000000000000000000000000000000001000000000000001000000000000000; // D (0x0000000040008000) 
    12'h332 : LOC <=          63'b000000000000000000000000000000001000000000000010000000000000000; // D (0x0000000040010000) 
    12'h471 : LOC <=          63'b000000000000000000000000000000001000000000000100000000000000000; // D (0x0000000040020000) 
    12'haf7 : LOC <=          63'b000000000000000000000000000000001000000000001000000000000000000; // D (0x0000000040040000) 
    12'h2c2 : LOC <=          63'b000000000000000000000000000000001000000000010000000000000000000; // D (0x0000000040080000) 
    12'h791 : LOC <=          63'b000000000000000000000000000000001000000000100000000000000000000; // D (0x0000000040100000) 
    12'hd37 : LOC <=          63'b000000000000000000000000000000001000000001000000000000000000000; // D (0x0000000040200000) 
    12'hd42 : LOC <=          63'b000000000000000000000000000000001000000010000000000000000000000; // D (0x0000000040400000) 
    12'hda8 : LOC <=          63'b000000000000000000000000000000001000000100000000000000000000000; // D (0x0000000040800000) 
    12'hc7c : LOC <=          63'b000000000000000000000000000000001000001000000000000000000000000; // D (0x0000000041000000) 
    12'hfd4 : LOC <=          63'b000000000000000000000000000000001000010000000000000000000000000; // D (0x0000000042000000) 
    12'h884 : LOC <=          63'b000000000000000000000000000000001000100000000000000000000000000; // D (0x0000000044000000) 
    12'h624 : LOC <=          63'b000000000000000000000000000000001001000000000000000000000000000; // D (0x0000000048000000) 
    12'he5d : LOC <=          63'b000000000000000000000000000000001010000000000000000000000000000; // D (0x0000000050000000) 
    12'hb96 : LOC <=          63'b000000000000000000000000000000001100000000000000000000000000000; // D (0x0000000060000000) 
    12'h1f3 : LOC <=          63'b000000000000000000000000000000001000000000000000000000000000000; // S (0x0000000040000000) 
//    12'h215 : LOC <=          63'b000000000000000000000000000000011000000000000000000000000000000; // D (0x00000000c0000000) 
//    12'h63f : LOC <=          63'b000000000000000000000000000000101000000000000000000000000000000; // D (0x0000000140000000) 
//    12'he6b : LOC <=          63'b000000000000000000000000000001001000000000000000000000000000000; // D (0x0000000240000000) 
//    12'hbfa : LOC <=          63'b000000000000000000000000000010001000000000000000000000000000000; // D (0x0000000440000000) 
//    12'h0d8 : LOC <=          63'b000000000000000000000000000100001000000000000000000000000000000; // D (0x0000000840000000) 
//    12'h3a5 : LOC <=          63'b000000000000000000000000001000001000000000000000000000000000000; // D (0x0000001040000000) 
//    12'h55f : LOC <=          63'b000000000000000000000000010000001000000000000000000000000000000; // D (0x0000002040000000) 
//    12'h8ab : LOC <=          63'b000000000000000000000000100000001000000000000000000000000000000; // D (0x0000004040000000) 
//    12'h67a : LOC <=          63'b000000000000000000000001000000001000000000000000000000000000000; // D (0x0000008040000000) 
//    12'hee1 : LOC <=          63'b000000000000000000000010000000001000000000000000000000000000000; // D (0x0000010040000000) 
//    12'haee : LOC <=          63'b000000000000000000000100000000001000000000000000000000000000000; // D (0x0000020040000000) 
//    12'h2f0 : LOC <=          63'b000000000000000000001000000000001000000000000000000000000000000; // D (0x0000040040000000) 
//    12'h7f5 : LOC <=          63'b000000000000000000010000000000001000000000000000000000000000000; // D (0x0000080040000000) 
//    12'hdff : LOC <=          63'b000000000000000000100000000000001000000000000000000000000000000; // D (0x0000100040000000) 
//    12'hcd2 : LOC <=          63'b000000000000000001000000000000001000000000000000000000000000000; // D (0x0000200040000000) 
//    12'he88 : LOC <=          63'b000000000000000010000000000000001000000000000000000000000000000; // D (0x0000400040000000) 
//    12'ha3c : LOC <=          63'b000000000000000100000000000000001000000000000000000000000000000; // D (0x0000800040000000) 
//    12'h354 : LOC <=          63'b000000000000001000000000000000001000000000000000000000000000000; // D (0x0001000040000000) 
//    12'h4bd : LOC <=          63'b000000000000010000000000000000001000000000000000000000000000000; // D (0x0002000040000000) 
//    12'hb6f : LOC <=          63'b000000000000100000000000000000001000000000000000000000000000000; // D (0x0004000040000000) 
//    12'h1f2 : LOC <=          63'b000000000001000000000000000000001000000000000000000000000000000; // D (0x0008000040000000) 
//    12'h1f1 : LOC <=          63'b000000000010000000000000000000001000000000000000000000000000000; // D (0x0010000040000000) 
//    12'h1f7 : LOC <=          63'b000000000100000000000000000000001000000000000000000000000000000; // D (0x0020000040000000) 
//    12'h1fb : LOC <=          63'b000000001000000000000000000000001000000000000000000000000000000; // D (0x0040000040000000) 
//    12'h1e3 : LOC <=          63'b000000010000000000000000000000001000000000000000000000000000000; // D (0x0080000040000000) 
//    12'h1d3 : LOC <=          63'b000000100000000000000000000000001000000000000000000000000000000; // D (0x0100000040000000) 
//    12'h1b3 : LOC <=          63'b000001000000000000000000000000001000000000000000000000000000000; // D (0x0200000040000000) 
//    12'h173 : LOC <=          63'b000010000000000000000000000000001000000000000000000000000000000; // D (0x0400000040000000) 
//    12'h0f3 : LOC <=          63'b000100000000000000000000000000001000000000000000000000000000000; // D (0x0800000040000000) 
//    12'h3f3 : LOC <=          63'b001000000000000000000000000000001000000000000000000000000000000; // D (0x1000000040000000) 
//    12'h5f3 : LOC <=          63'b010000000000000000000000000000001000000000000000000000000000000; // D (0x2000000040000000) 
//    12'h9f3 : LOC <=          63'b100000000000000000000000000000001000000000000000000000000000000; // D (0x4000000040000000) 
    12'h6df : LOC <=          63'b000000000000000000000000000000010000000000000000000000000000001; // D (0x0000000080000001) 
    12'h994 : LOC <=          63'b000000000000000000000000000000010000000000000000000000000000010; // D (0x0000000080000002) 
    12'h23b : LOC <=          63'b000000000000000000000000000000010000000000000000000000000000100; // D (0x0000000080000004) 
    12'h05c : LOC <=          63'b000000000000000000000000000000010000000000000000000000000001000; // D (0x0000000080000008) 
    12'h492 : LOC <=          63'b000000000000000000000000000000010000000000000000000000000010000; // D (0x0000000080000010) 
    12'hd0e : LOC <=          63'b000000000000000000000000000000010000000000000000000000000100000; // D (0x0000000080000020) 
    12'hb0f : LOC <=          63'b000000000000000000000000000000010000000000000000000000001000000; // D (0x0000000080000040) 
    12'h70d : LOC <=          63'b000000000000000000000000000000010000000000000000000000010000000; // D (0x0000000080000080) 
    12'ha30 : LOC <=          63'b000000000000000000000000000000010000000000000000000000100000000; // D (0x0000000080000100) 
    12'h573 : LOC <=          63'b000000000000000000000000000000010000000000000000000001000000000; // D (0x0000000080000200) 
    12'hecc : LOC <=          63'b000000000000000000000000000000010000000000000000000010000000000; // D (0x0000000080000400) 
    12'hc8b : LOC <=          63'b000000000000000000000000000000010000000000000000000100000000000; // D (0x0000000080000800) 
    12'h805 : LOC <=          63'b000000000000000000000000000000010000000000000000001000000000000; // D (0x0000000080001000) 
    12'h119 : LOC <=          63'b000000000000000000000000000000010000000000000000010000000000000; // D (0x0000000080002000) 
    12'h618 : LOC <=          63'b000000000000000000000000000000010000000000000000100000000000000; // D (0x0000000080004000) 
    12'h81a : LOC <=          63'b000000000000000000000000000000010000000000000001000000000000000; // D (0x0000000080008000) 
    12'h127 : LOC <=          63'b000000000000000000000000000000010000000000000010000000000000000; // D (0x0000000080010000) 
    12'h664 : LOC <=          63'b000000000000000000000000000000010000000000000100000000000000000; // D (0x0000000080020000) 
    12'h8e2 : LOC <=          63'b000000000000000000000000000000010000000000001000000000000000000; // D (0x0000000080040000) 
    12'h0d7 : LOC <=          63'b000000000000000000000000000000010000000000010000000000000000000; // D (0x0000000080080000) 
    12'h584 : LOC <=          63'b000000000000000000000000000000010000000000100000000000000000000; // D (0x0000000080100000) 
    12'hf22 : LOC <=          63'b000000000000000000000000000000010000000001000000000000000000000; // D (0x0000000080200000) 
    12'hf57 : LOC <=          63'b000000000000000000000000000000010000000010000000000000000000000; // D (0x0000000080400000) 
    12'hfbd : LOC <=          63'b000000000000000000000000000000010000000100000000000000000000000; // D (0x0000000080800000) 
    12'he69 : LOC <=          63'b000000000000000000000000000000010000001000000000000000000000000; // D (0x0000000081000000) 
    12'hdc1 : LOC <=          63'b000000000000000000000000000000010000010000000000000000000000000; // D (0x0000000082000000) 
    12'ha91 : LOC <=          63'b000000000000000000000000000000010000100000000000000000000000000; // D (0x0000000084000000) 
    12'h431 : LOC <=          63'b000000000000000000000000000000010001000000000000000000000000000; // D (0x0000000088000000) 
    12'hc48 : LOC <=          63'b000000000000000000000000000000010010000000000000000000000000000; // D (0x0000000090000000) 
    12'h983 : LOC <=          63'b000000000000000000000000000000010100000000000000000000000000000; // D (0x00000000a0000000) 
    12'h215 : LOC <=          63'b000000000000000000000000000000011000000000000000000000000000000; // D (0x00000000c0000000) 
    12'h3e6 : LOC <=          63'b000000000000000000000000000000010000000000000000000000000000000; // S (0x0000000080000000) 
//    12'h42a : LOC <=          63'b000000000000000000000000000000110000000000000000000000000000000; // D (0x0000000180000000) 
//    12'hc7e : LOC <=          63'b000000000000000000000000000001010000000000000000000000000000000; // D (0x0000000280000000) 
//    12'h9ef : LOC <=          63'b000000000000000000000000000010010000000000000000000000000000000; // D (0x0000000480000000) 
//    12'h2cd : LOC <=          63'b000000000000000000000000000100010000000000000000000000000000000; // D (0x0000000880000000) 
//    12'h1b0 : LOC <=          63'b000000000000000000000000001000010000000000000000000000000000000; // D (0x0000001080000000) 
//    12'h74a : LOC <=          63'b000000000000000000000000010000010000000000000000000000000000000; // D (0x0000002080000000) 
//    12'habe : LOC <=          63'b000000000000000000000000100000010000000000000000000000000000000; // D (0x0000004080000000) 
//    12'h46f : LOC <=          63'b000000000000000000000001000000010000000000000000000000000000000; // D (0x0000008080000000) 
//    12'hcf4 : LOC <=          63'b000000000000000000000010000000010000000000000000000000000000000; // D (0x0000010080000000) 
//    12'h8fb : LOC <=          63'b000000000000000000000100000000010000000000000000000000000000000; // D (0x0000020080000000) 
//    12'h0e5 : LOC <=          63'b000000000000000000001000000000010000000000000000000000000000000; // D (0x0000040080000000) 
//    12'h5e0 : LOC <=          63'b000000000000000000010000000000010000000000000000000000000000000; // D (0x0000080080000000) 
//    12'hfea : LOC <=          63'b000000000000000000100000000000010000000000000000000000000000000; // D (0x0000100080000000) 
//    12'hec7 : LOC <=          63'b000000000000000001000000000000010000000000000000000000000000000; // D (0x0000200080000000) 
//    12'hc9d : LOC <=          63'b000000000000000010000000000000010000000000000000000000000000000; // D (0x0000400080000000) 
//    12'h829 : LOC <=          63'b000000000000000100000000000000010000000000000000000000000000000; // D (0x0000800080000000) 
//    12'h141 : LOC <=          63'b000000000000001000000000000000010000000000000000000000000000000; // D (0x0001000080000000) 
//    12'h6a8 : LOC <=          63'b000000000000010000000000000000010000000000000000000000000000000; // D (0x0002000080000000) 
//    12'h97a : LOC <=          63'b000000000000100000000000000000010000000000000000000000000000000; // D (0x0004000080000000) 
//    12'h3e7 : LOC <=          63'b000000000001000000000000000000010000000000000000000000000000000; // D (0x0008000080000000) 
//    12'h3e4 : LOC <=          63'b000000000010000000000000000000010000000000000000000000000000000; // D (0x0010000080000000) 
//    12'h3e2 : LOC <=          63'b000000000100000000000000000000010000000000000000000000000000000; // D (0x0020000080000000) 
//    12'h3ee : LOC <=          63'b000000001000000000000000000000010000000000000000000000000000000; // D (0x0040000080000000) 
//    12'h3f6 : LOC <=          63'b000000010000000000000000000000010000000000000000000000000000000; // D (0x0080000080000000) 
//    12'h3c6 : LOC <=          63'b000000100000000000000000000000010000000000000000000000000000000; // D (0x0100000080000000) 
//    12'h3a6 : LOC <=          63'b000001000000000000000000000000010000000000000000000000000000000; // D (0x0200000080000000) 
//    12'h366 : LOC <=          63'b000010000000000000000000000000010000000000000000000000000000000; // D (0x0400000080000000) 
//    12'h2e6 : LOC <=          63'b000100000000000000000000000000010000000000000000000000000000000; // D (0x0800000080000000) 
//    12'h1e6 : LOC <=          63'b001000000000000000000000000000010000000000000000000000000000000; // D (0x1000000080000000) 
//    12'h7e6 : LOC <=          63'b010000000000000000000000000000010000000000000000000000000000000; // D (0x2000000080000000) 
//    12'hbe6 : LOC <=          63'b100000000000000000000000000000010000000000000000000000000000000; // D (0x4000000080000000) 
    12'h2f5 : LOC <=          63'b000000000000000000000000000000100000000000000000000000000000001; // D (0x0000000100000001) 
    12'hdbe : LOC <=          63'b000000000000000000000000000000100000000000000000000000000000010; // D (0x0000000100000002) 
    12'h611 : LOC <=          63'b000000000000000000000000000000100000000000000000000000000000100; // D (0x0000000100000004) 
    12'h476 : LOC <=          63'b000000000000000000000000000000100000000000000000000000000001000; // D (0x0000000100000008) 
    12'h0b8 : LOC <=          63'b000000000000000000000000000000100000000000000000000000000010000; // D (0x0000000100000010) 
    12'h924 : LOC <=          63'b000000000000000000000000000000100000000000000000000000000100000; // D (0x0000000100000020) 
    12'hf25 : LOC <=          63'b000000000000000000000000000000100000000000000000000000001000000; // D (0x0000000100000040) 
    12'h327 : LOC <=          63'b000000000000000000000000000000100000000000000000000000010000000; // D (0x0000000100000080) 
    12'he1a : LOC <=          63'b000000000000000000000000000000100000000000000000000000100000000; // D (0x0000000100000100) 
    12'h159 : LOC <=          63'b000000000000000000000000000000100000000000000000000001000000000; // D (0x0000000100000200) 
    12'hae6 : LOC <=          63'b000000000000000000000000000000100000000000000000000010000000000; // D (0x0000000100000400) 
    12'h8a1 : LOC <=          63'b000000000000000000000000000000100000000000000000000100000000000; // D (0x0000000100000800) 
    12'hc2f : LOC <=          63'b000000000000000000000000000000100000000000000000001000000000000; // D (0x0000000100001000) 
    12'h533 : LOC <=          63'b000000000000000000000000000000100000000000000000010000000000000; // D (0x0000000100002000) 
    12'h232 : LOC <=          63'b000000000000000000000000000000100000000000000000100000000000000; // D (0x0000000100004000) 
    12'hc30 : LOC <=          63'b000000000000000000000000000000100000000000000001000000000000000; // D (0x0000000100008000) 
    12'h50d : LOC <=          63'b000000000000000000000000000000100000000000000010000000000000000; // D (0x0000000100010000) 
    12'h24e : LOC <=          63'b000000000000000000000000000000100000000000000100000000000000000; // D (0x0000000100020000) 
    12'hcc8 : LOC <=          63'b000000000000000000000000000000100000000000001000000000000000000; // D (0x0000000100040000) 
    12'h4fd : LOC <=          63'b000000000000000000000000000000100000000000010000000000000000000; // D (0x0000000100080000) 
    12'h1ae : LOC <=          63'b000000000000000000000000000000100000000000100000000000000000000; // D (0x0000000100100000) 
    12'hb08 : LOC <=          63'b000000000000000000000000000000100000000001000000000000000000000; // D (0x0000000100200000) 
    12'hb7d : LOC <=          63'b000000000000000000000000000000100000000010000000000000000000000; // D (0x0000000100400000) 
    12'hb97 : LOC <=          63'b000000000000000000000000000000100000000100000000000000000000000; // D (0x0000000100800000) 
    12'ha43 : LOC <=          63'b000000000000000000000000000000100000001000000000000000000000000; // D (0x0000000101000000) 
    12'h9eb : LOC <=          63'b000000000000000000000000000000100000010000000000000000000000000; // D (0x0000000102000000) 
    12'hebb : LOC <=          63'b000000000000000000000000000000100000100000000000000000000000000; // D (0x0000000104000000) 
    12'h01b : LOC <=          63'b000000000000000000000000000000100001000000000000000000000000000; // D (0x0000000108000000) 
    12'h862 : LOC <=          63'b000000000000000000000000000000100010000000000000000000000000000; // D (0x0000000110000000) 
    12'hda9 : LOC <=          63'b000000000000000000000000000000100100000000000000000000000000000; // D (0x0000000120000000) 
    12'h63f : LOC <=          63'b000000000000000000000000000000101000000000000000000000000000000; // D (0x0000000140000000) 
    12'h42a : LOC <=          63'b000000000000000000000000000000110000000000000000000000000000000; // D (0x0000000180000000) 
    12'h7cc : LOC <=          63'b000000000000000000000000000000100000000000000000000000000000000; // S (0x0000000100000000) 
//    12'h854 : LOC <=          63'b000000000000000000000000000001100000000000000000000000000000000; // D (0x0000000300000000) 
//    12'hdc5 : LOC <=          63'b000000000000000000000000000010100000000000000000000000000000000; // D (0x0000000500000000) 
//    12'h6e7 : LOC <=          63'b000000000000000000000000000100100000000000000000000000000000000; // D (0x0000000900000000) 
//    12'h59a : LOC <=          63'b000000000000000000000000001000100000000000000000000000000000000; // D (0x0000001100000000) 
//    12'h360 : LOC <=          63'b000000000000000000000000010000100000000000000000000000000000000; // D (0x0000002100000000) 
//    12'he94 : LOC <=          63'b000000000000000000000000100000100000000000000000000000000000000; // D (0x0000004100000000) 
//    12'h045 : LOC <=          63'b000000000000000000000001000000100000000000000000000000000000000; // D (0x0000008100000000) 
//    12'h8de : LOC <=          63'b000000000000000000000010000000100000000000000000000000000000000; // D (0x0000010100000000) 
//    12'hcd1 : LOC <=          63'b000000000000000000000100000000100000000000000000000000000000000; // D (0x0000020100000000) 
//    12'h4cf : LOC <=          63'b000000000000000000001000000000100000000000000000000000000000000; // D (0x0000040100000000) 
//    12'h1ca : LOC <=          63'b000000000000000000010000000000100000000000000000000000000000000; // D (0x0000080100000000) 
//    12'hbc0 : LOC <=          63'b000000000000000000100000000000100000000000000000000000000000000; // D (0x0000100100000000) 
//    12'haed : LOC <=          63'b000000000000000001000000000000100000000000000000000000000000000; // D (0x0000200100000000) 
//    12'h8b7 : LOC <=          63'b000000000000000010000000000000100000000000000000000000000000000; // D (0x0000400100000000) 
//    12'hc03 : LOC <=          63'b000000000000000100000000000000100000000000000000000000000000000; // D (0x0000800100000000) 
//    12'h56b : LOC <=          63'b000000000000001000000000000000100000000000000000000000000000000; // D (0x0001000100000000) 
//    12'h282 : LOC <=          63'b000000000000010000000000000000100000000000000000000000000000000; // D (0x0002000100000000) 
//    12'hd50 : LOC <=          63'b000000000000100000000000000000100000000000000000000000000000000; // D (0x0004000100000000) 
//    12'h7cd : LOC <=          63'b000000000001000000000000000000100000000000000000000000000000000; // D (0x0008000100000000) 
//    12'h7ce : LOC <=          63'b000000000010000000000000000000100000000000000000000000000000000; // D (0x0010000100000000) 
//    12'h7c8 : LOC <=          63'b000000000100000000000000000000100000000000000000000000000000000; // D (0x0020000100000000) 
//    12'h7c4 : LOC <=          63'b000000001000000000000000000000100000000000000000000000000000000; // D (0x0040000100000000) 
//    12'h7dc : LOC <=          63'b000000010000000000000000000000100000000000000000000000000000000; // D (0x0080000100000000) 
//    12'h7ec : LOC <=          63'b000000100000000000000000000000100000000000000000000000000000000; // D (0x0100000100000000) 
//    12'h78c : LOC <=          63'b000001000000000000000000000000100000000000000000000000000000000; // D (0x0200000100000000) 
//    12'h74c : LOC <=          63'b000010000000000000000000000000100000000000000000000000000000000; // D (0x0400000100000000) 
//    12'h6cc : LOC <=          63'b000100000000000000000000000000100000000000000000000000000000000; // D (0x0800000100000000) 
//    12'h5cc : LOC <=          63'b001000000000000000000000000000100000000000000000000000000000000; // D (0x1000000100000000) 
//    12'h3cc : LOC <=          63'b010000000000000000000000000000100000000000000000000000000000000; // D (0x2000000100000000) 
//    12'hfcc : LOC <=          63'b100000000000000000000000000000100000000000000000000000000000000; // D (0x4000000100000000) 
    12'haa1 : LOC <=          63'b000000000000000000000000000001000000000000000000000000000000001; // D (0x0000000200000001) 
    12'h5ea : LOC <=          63'b000000000000000000000000000001000000000000000000000000000000010; // D (0x0000000200000002) 
    12'he45 : LOC <=          63'b000000000000000000000000000001000000000000000000000000000000100; // D (0x0000000200000004) 
    12'hc22 : LOC <=          63'b000000000000000000000000000001000000000000000000000000000001000; // D (0x0000000200000008) 
    12'h8ec : LOC <=          63'b000000000000000000000000000001000000000000000000000000000010000; // D (0x0000000200000010) 
    12'h170 : LOC <=          63'b000000000000000000000000000001000000000000000000000000000100000; // D (0x0000000200000020) 
    12'h771 : LOC <=          63'b000000000000000000000000000001000000000000000000000000001000000; // D (0x0000000200000040) 
    12'hb73 : LOC <=          63'b000000000000000000000000000001000000000000000000000000010000000; // D (0x0000000200000080) 
    12'h64e : LOC <=          63'b000000000000000000000000000001000000000000000000000000100000000; // D (0x0000000200000100) 
    12'h90d : LOC <=          63'b000000000000000000000000000001000000000000000000000001000000000; // D (0x0000000200000200) 
    12'h2b2 : LOC <=          63'b000000000000000000000000000001000000000000000000000010000000000; // D (0x0000000200000400) 
    12'h0f5 : LOC <=          63'b000000000000000000000000000001000000000000000000000100000000000; // D (0x0000000200000800) 
    12'h47b : LOC <=          63'b000000000000000000000000000001000000000000000000001000000000000; // D (0x0000000200001000) 
    12'hd67 : LOC <=          63'b000000000000000000000000000001000000000000000000010000000000000; // D (0x0000000200002000) 
    12'ha66 : LOC <=          63'b000000000000000000000000000001000000000000000000100000000000000; // D (0x0000000200004000) 
    12'h464 : LOC <=          63'b000000000000000000000000000001000000000000000001000000000000000; // D (0x0000000200008000) 
    12'hd59 : LOC <=          63'b000000000000000000000000000001000000000000000010000000000000000; // D (0x0000000200010000) 
    12'ha1a : LOC <=          63'b000000000000000000000000000001000000000000000100000000000000000; // D (0x0000000200020000) 
    12'h49c : LOC <=          63'b000000000000000000000000000001000000000000001000000000000000000; // D (0x0000000200040000) 
    12'hca9 : LOC <=          63'b000000000000000000000000000001000000000000010000000000000000000; // D (0x0000000200080000) 
    12'h9fa : LOC <=          63'b000000000000000000000000000001000000000000100000000000000000000; // D (0x0000000200100000) 
    12'h35c : LOC <=          63'b000000000000000000000000000001000000000001000000000000000000000; // D (0x0000000200200000) 
    12'h329 : LOC <=          63'b000000000000000000000000000001000000000010000000000000000000000; // D (0x0000000200400000) 
    12'h3c3 : LOC <=          63'b000000000000000000000000000001000000000100000000000000000000000; // D (0x0000000200800000) 
    12'h217 : LOC <=          63'b000000000000000000000000000001000000001000000000000000000000000; // D (0x0000000201000000) 
    12'h1bf : LOC <=          63'b000000000000000000000000000001000000010000000000000000000000000; // D (0x0000000202000000) 
    12'h6ef : LOC <=          63'b000000000000000000000000000001000000100000000000000000000000000; // D (0x0000000204000000) 
    12'h84f : LOC <=          63'b000000000000000000000000000001000001000000000000000000000000000; // D (0x0000000208000000) 
    12'h036 : LOC <=          63'b000000000000000000000000000001000010000000000000000000000000000; // D (0x0000000210000000) 
    12'h5fd : LOC <=          63'b000000000000000000000000000001000100000000000000000000000000000; // D (0x0000000220000000) 
    12'he6b : LOC <=          63'b000000000000000000000000000001001000000000000000000000000000000; // D (0x0000000240000000) 
    12'hc7e : LOC <=          63'b000000000000000000000000000001010000000000000000000000000000000; // D (0x0000000280000000) 
    12'h854 : LOC <=          63'b000000000000000000000000000001100000000000000000000000000000000; // D (0x0000000300000000) 
    12'hf98 : LOC <=          63'b000000000000000000000000000001000000000000000000000000000000000; // S (0x0000000200000000) 
//    12'h591 : LOC <=          63'b000000000000000000000000000011000000000000000000000000000000000; // D (0x0000000600000000) 
//    12'heb3 : LOC <=          63'b000000000000000000000000000101000000000000000000000000000000000; // D (0x0000000a00000000) 
//    12'hdce : LOC <=          63'b000000000000000000000000001001000000000000000000000000000000000; // D (0x0000001200000000) 
//    12'hb34 : LOC <=          63'b000000000000000000000000010001000000000000000000000000000000000; // D (0x0000002200000000) 
//    12'h6c0 : LOC <=          63'b000000000000000000000000100001000000000000000000000000000000000; // D (0x0000004200000000) 
//    12'h811 : LOC <=          63'b000000000000000000000001000001000000000000000000000000000000000; // D (0x0000008200000000) 
//    12'h08a : LOC <=          63'b000000000000000000000010000001000000000000000000000000000000000; // D (0x0000010200000000) 
//    12'h485 : LOC <=          63'b000000000000000000000100000001000000000000000000000000000000000; // D (0x0000020200000000) 
//    12'hc9b : LOC <=          63'b000000000000000000001000000001000000000000000000000000000000000; // D (0x0000040200000000) 
//    12'h99e : LOC <=          63'b000000000000000000010000000001000000000000000000000000000000000; // D (0x0000080200000000) 
//    12'h394 : LOC <=          63'b000000000000000000100000000001000000000000000000000000000000000; // D (0x0000100200000000) 
//    12'h2b9 : LOC <=          63'b000000000000000001000000000001000000000000000000000000000000000; // D (0x0000200200000000) 
//    12'h0e3 : LOC <=          63'b000000000000000010000000000001000000000000000000000000000000000; // D (0x0000400200000000) 
//    12'h457 : LOC <=          63'b000000000000000100000000000001000000000000000000000000000000000; // D (0x0000800200000000) 
//    12'hd3f : LOC <=          63'b000000000000001000000000000001000000000000000000000000000000000; // D (0x0001000200000000) 
//    12'had6 : LOC <=          63'b000000000000010000000000000001000000000000000000000000000000000; // D (0x0002000200000000) 
//    12'h504 : LOC <=          63'b000000000000100000000000000001000000000000000000000000000000000; // D (0x0004000200000000) 
//    12'hf99 : LOC <=          63'b000000000001000000000000000001000000000000000000000000000000000; // D (0x0008000200000000) 
//    12'hf9a : LOC <=          63'b000000000010000000000000000001000000000000000000000000000000000; // D (0x0010000200000000) 
//    12'hf9c : LOC <=          63'b000000000100000000000000000001000000000000000000000000000000000; // D (0x0020000200000000) 
//    12'hf90 : LOC <=          63'b000000001000000000000000000001000000000000000000000000000000000; // D (0x0040000200000000) 
//    12'hf88 : LOC <=          63'b000000010000000000000000000001000000000000000000000000000000000; // D (0x0080000200000000) 
//    12'hfb8 : LOC <=          63'b000000100000000000000000000001000000000000000000000000000000000; // D (0x0100000200000000) 
//    12'hfd8 : LOC <=          63'b000001000000000000000000000001000000000000000000000000000000000; // D (0x0200000200000000) 
//    12'hf18 : LOC <=          63'b000010000000000000000000000001000000000000000000000000000000000; // D (0x0400000200000000) 
//    12'he98 : LOC <=          63'b000100000000000000000000000001000000000000000000000000000000000; // D (0x0800000200000000) 
//    12'hd98 : LOC <=          63'b001000000000000000000000000001000000000000000000000000000000000; // D (0x1000000200000000) 
//    12'hb98 : LOC <=          63'b010000000000000000000000000001000000000000000000000000000000000; // D (0x2000000200000000) 
//    12'h798 : LOC <=          63'b100000000000000000000000000001000000000000000000000000000000000; // D (0x4000000200000000) 
    12'hf30 : LOC <=          63'b000000000000000000000000000010000000000000000000000000000000001; // D (0x0000000400000001) 
    12'h07b : LOC <=          63'b000000000000000000000000000010000000000000000000000000000000010; // D (0x0000000400000002) 
    12'hbd4 : LOC <=          63'b000000000000000000000000000010000000000000000000000000000000100; // D (0x0000000400000004) 
    12'h9b3 : LOC <=          63'b000000000000000000000000000010000000000000000000000000000001000; // D (0x0000000400000008) 
    12'hd7d : LOC <=          63'b000000000000000000000000000010000000000000000000000000000010000; // D (0x0000000400000010) 
    12'h4e1 : LOC <=          63'b000000000000000000000000000010000000000000000000000000000100000; // D (0x0000000400000020) 
    12'h2e0 : LOC <=          63'b000000000000000000000000000010000000000000000000000000001000000; // D (0x0000000400000040) 
    12'hee2 : LOC <=          63'b000000000000000000000000000010000000000000000000000000010000000; // D (0x0000000400000080) 
    12'h3df : LOC <=          63'b000000000000000000000000000010000000000000000000000000100000000; // D (0x0000000400000100) 
    12'hc9c : LOC <=          63'b000000000000000000000000000010000000000000000000000001000000000; // D (0x0000000400000200) 
    12'h723 : LOC <=          63'b000000000000000000000000000010000000000000000000000010000000000; // D (0x0000000400000400) 
    12'h564 : LOC <=          63'b000000000000000000000000000010000000000000000000000100000000000; // D (0x0000000400000800) 
    12'h1ea : LOC <=          63'b000000000000000000000000000010000000000000000000001000000000000; // D (0x0000000400001000) 
    12'h8f6 : LOC <=          63'b000000000000000000000000000010000000000000000000010000000000000; // D (0x0000000400002000) 
    12'hff7 : LOC <=          63'b000000000000000000000000000010000000000000000000100000000000000; // D (0x0000000400004000) 
    12'h1f5 : LOC <=          63'b000000000000000000000000000010000000000000000001000000000000000; // D (0x0000000400008000) 
    12'h8c8 : LOC <=          63'b000000000000000000000000000010000000000000000010000000000000000; // D (0x0000000400010000) 
    12'hf8b : LOC <=          63'b000000000000000000000000000010000000000000000100000000000000000; // D (0x0000000400020000) 
    12'h10d : LOC <=          63'b000000000000000000000000000010000000000000001000000000000000000; // D (0x0000000400040000) 
    12'h938 : LOC <=          63'b000000000000000000000000000010000000000000010000000000000000000; // D (0x0000000400080000) 
    12'hc6b : LOC <=          63'b000000000000000000000000000010000000000000100000000000000000000; // D (0x0000000400100000) 
    12'h6cd : LOC <=          63'b000000000000000000000000000010000000000001000000000000000000000; // D (0x0000000400200000) 
    12'h6b8 : LOC <=          63'b000000000000000000000000000010000000000010000000000000000000000; // D (0x0000000400400000) 
    12'h652 : LOC <=          63'b000000000000000000000000000010000000000100000000000000000000000; // D (0x0000000400800000) 
    12'h786 : LOC <=          63'b000000000000000000000000000010000000001000000000000000000000000; // D (0x0000000401000000) 
    12'h42e : LOC <=          63'b000000000000000000000000000010000000010000000000000000000000000; // D (0x0000000402000000) 
    12'h37e : LOC <=          63'b000000000000000000000000000010000000100000000000000000000000000; // D (0x0000000404000000) 
    12'hdde : LOC <=          63'b000000000000000000000000000010000001000000000000000000000000000; // D (0x0000000408000000) 
    12'h5a7 : LOC <=          63'b000000000000000000000000000010000010000000000000000000000000000; // D (0x0000000410000000) 
    12'h06c : LOC <=          63'b000000000000000000000000000010000100000000000000000000000000000; // D (0x0000000420000000) 
    12'hbfa : LOC <=          63'b000000000000000000000000000010001000000000000000000000000000000; // D (0x0000000440000000) 
    12'h9ef : LOC <=          63'b000000000000000000000000000010010000000000000000000000000000000; // D (0x0000000480000000) 
    12'hdc5 : LOC <=          63'b000000000000000000000000000010100000000000000000000000000000000; // D (0x0000000500000000) 
    12'h591 : LOC <=          63'b000000000000000000000000000011000000000000000000000000000000000; // D (0x0000000600000000) 
    12'ha09 : LOC <=          63'b000000000000000000000000000010000000000000000000000000000000000; // S (0x0000000400000000) 
//    12'hb22 : LOC <=          63'b000000000000000000000000000110000000000000000000000000000000000; // D (0x0000000c00000000) 
//    12'h85f : LOC <=          63'b000000000000000000000000001010000000000000000000000000000000000; // D (0x0000001400000000) 
//    12'hea5 : LOC <=          63'b000000000000000000000000010010000000000000000000000000000000000; // D (0x0000002400000000) 
//    12'h351 : LOC <=          63'b000000000000000000000000100010000000000000000000000000000000000; // D (0x0000004400000000) 
//    12'hd80 : LOC <=          63'b000000000000000000000001000010000000000000000000000000000000000; // D (0x0000008400000000) 
//    12'h51b : LOC <=          63'b000000000000000000000010000010000000000000000000000000000000000; // D (0x0000010400000000) 
//    12'h114 : LOC <=          63'b000000000000000000000100000010000000000000000000000000000000000; // D (0x0000020400000000) 
//    12'h90a : LOC <=          63'b000000000000000000001000000010000000000000000000000000000000000; // D (0x0000040400000000) 
//    12'hc0f : LOC <=          63'b000000000000000000010000000010000000000000000000000000000000000; // D (0x0000080400000000) 
//    12'h605 : LOC <=          63'b000000000000000000100000000010000000000000000000000000000000000; // D (0x0000100400000000) 
//    12'h728 : LOC <=          63'b000000000000000001000000000010000000000000000000000000000000000; // D (0x0000200400000000) 
//    12'h572 : LOC <=          63'b000000000000000010000000000010000000000000000000000000000000000; // D (0x0000400400000000) 
//    12'h1c6 : LOC <=          63'b000000000000000100000000000010000000000000000000000000000000000; // D (0x0000800400000000) 
//    12'h8ae : LOC <=          63'b000000000000001000000000000010000000000000000000000000000000000; // D (0x0001000400000000) 
//    12'hf47 : LOC <=          63'b000000000000010000000000000010000000000000000000000000000000000; // D (0x0002000400000000) 
//    12'h095 : LOC <=          63'b000000000000100000000000000010000000000000000000000000000000000; // D (0x0004000400000000) 
//    12'ha08 : LOC <=          63'b000000000001000000000000000010000000000000000000000000000000000; // D (0x0008000400000000) 
//    12'ha0b : LOC <=          63'b000000000010000000000000000010000000000000000000000000000000000; // D (0x0010000400000000) 
//    12'ha0d : LOC <=          63'b000000000100000000000000000010000000000000000000000000000000000; // D (0x0020000400000000) 
//    12'ha01 : LOC <=          63'b000000001000000000000000000010000000000000000000000000000000000; // D (0x0040000400000000) 
//    12'ha19 : LOC <=          63'b000000010000000000000000000010000000000000000000000000000000000; // D (0x0080000400000000) 
//    12'ha29 : LOC <=          63'b000000100000000000000000000010000000000000000000000000000000000; // D (0x0100000400000000) 
//    12'ha49 : LOC <=          63'b000001000000000000000000000010000000000000000000000000000000000; // D (0x0200000400000000) 
//    12'ha89 : LOC <=          63'b000010000000000000000000000010000000000000000000000000000000000; // D (0x0400000400000000) 
//    12'hb09 : LOC <=          63'b000100000000000000000000000010000000000000000000000000000000000; // D (0x0800000400000000) 
//    12'h809 : LOC <=          63'b001000000000000000000000000010000000000000000000000000000000000; // D (0x1000000400000000) 
//    12'he09 : LOC <=          63'b010000000000000000000000000010000000000000000000000000000000000; // D (0x2000000400000000) 
//    12'h209 : LOC <=          63'b100000000000000000000000000010000000000000000000000000000000000; // D (0x4000000400000000) 
    12'h412 : LOC <=          63'b000000000000000000000000000100000000000000000000000000000000001; // D (0x0000000800000001) 
    12'hb59 : LOC <=          63'b000000000000000000000000000100000000000000000000000000000000010; // D (0x0000000800000002) 
    12'h0f6 : LOC <=          63'b000000000000000000000000000100000000000000000000000000000000100; // D (0x0000000800000004) 
    12'h291 : LOC <=          63'b000000000000000000000000000100000000000000000000000000000001000; // D (0x0000000800000008) 
    12'h65f : LOC <=          63'b000000000000000000000000000100000000000000000000000000000010000; // D (0x0000000800000010) 
    12'hfc3 : LOC <=          63'b000000000000000000000000000100000000000000000000000000000100000; // D (0x0000000800000020) 
    12'h9c2 : LOC <=          63'b000000000000000000000000000100000000000000000000000000001000000; // D (0x0000000800000040) 
    12'h5c0 : LOC <=          63'b000000000000000000000000000100000000000000000000000000010000000; // D (0x0000000800000080) 
    12'h8fd : LOC <=          63'b000000000000000000000000000100000000000000000000000000100000000; // D (0x0000000800000100) 
    12'h7be : LOC <=          63'b000000000000000000000000000100000000000000000000000001000000000; // D (0x0000000800000200) 
    12'hc01 : LOC <=          63'b000000000000000000000000000100000000000000000000000010000000000; // D (0x0000000800000400) 
    12'he46 : LOC <=          63'b000000000000000000000000000100000000000000000000000100000000000; // D (0x0000000800000800) 
    12'hac8 : LOC <=          63'b000000000000000000000000000100000000000000000000001000000000000; // D (0x0000000800001000) 
    12'h3d4 : LOC <=          63'b000000000000000000000000000100000000000000000000010000000000000; // D (0x0000000800002000) 
    12'h4d5 : LOC <=          63'b000000000000000000000000000100000000000000000000100000000000000; // D (0x0000000800004000) 
    12'had7 : LOC <=          63'b000000000000000000000000000100000000000000000001000000000000000; // D (0x0000000800008000) 
    12'h3ea : LOC <=          63'b000000000000000000000000000100000000000000000010000000000000000; // D (0x0000000800010000) 
    12'h4a9 : LOC <=          63'b000000000000000000000000000100000000000000000100000000000000000; // D (0x0000000800020000) 
    12'ha2f : LOC <=          63'b000000000000000000000000000100000000000000001000000000000000000; // D (0x0000000800040000) 
    12'h21a : LOC <=          63'b000000000000000000000000000100000000000000010000000000000000000; // D (0x0000000800080000) 
    12'h749 : LOC <=          63'b000000000000000000000000000100000000000000100000000000000000000; // D (0x0000000800100000) 
    12'hdef : LOC <=          63'b000000000000000000000000000100000000000001000000000000000000000; // D (0x0000000800200000) 
    12'hd9a : LOC <=          63'b000000000000000000000000000100000000000010000000000000000000000; // D (0x0000000800400000) 
    12'hd70 : LOC <=          63'b000000000000000000000000000100000000000100000000000000000000000; // D (0x0000000800800000) 
    12'hca4 : LOC <=          63'b000000000000000000000000000100000000001000000000000000000000000; // D (0x0000000801000000) 
    12'hf0c : LOC <=          63'b000000000000000000000000000100000000010000000000000000000000000; // D (0x0000000802000000) 
    12'h85c : LOC <=          63'b000000000000000000000000000100000000100000000000000000000000000; // D (0x0000000804000000) 
    12'h6fc : LOC <=          63'b000000000000000000000000000100000001000000000000000000000000000; // D (0x0000000808000000) 
    12'he85 : LOC <=          63'b000000000000000000000000000100000010000000000000000000000000000; // D (0x0000000810000000) 
    12'hb4e : LOC <=          63'b000000000000000000000000000100000100000000000000000000000000000; // D (0x0000000820000000) 
    12'h0d8 : LOC <=          63'b000000000000000000000000000100001000000000000000000000000000000; // D (0x0000000840000000) 
    12'h2cd : LOC <=          63'b000000000000000000000000000100010000000000000000000000000000000; // D (0x0000000880000000) 
    12'h6e7 : LOC <=          63'b000000000000000000000000000100100000000000000000000000000000000; // D (0x0000000900000000) 
    12'heb3 : LOC <=          63'b000000000000000000000000000101000000000000000000000000000000000; // D (0x0000000a00000000) 
    12'hb22 : LOC <=          63'b000000000000000000000000000110000000000000000000000000000000000; // D (0x0000000c00000000) 
    12'h12b : LOC <=          63'b000000000000000000000000000100000000000000000000000000000000000; // S (0x0000000800000000) 
//    12'h37d : LOC <=          63'b000000000000000000000000001100000000000000000000000000000000000; // D (0x0000001800000000) 
//    12'h587 : LOC <=          63'b000000000000000000000000010100000000000000000000000000000000000; // D (0x0000002800000000) 
//    12'h873 : LOC <=          63'b000000000000000000000000100100000000000000000000000000000000000; // D (0x0000004800000000) 
//    12'h6a2 : LOC <=          63'b000000000000000000000001000100000000000000000000000000000000000; // D (0x0000008800000000) 
//    12'he39 : LOC <=          63'b000000000000000000000010000100000000000000000000000000000000000; // D (0x0000010800000000) 
//    12'ha36 : LOC <=          63'b000000000000000000000100000100000000000000000000000000000000000; // D (0x0000020800000000) 
//    12'h228 : LOC <=          63'b000000000000000000001000000100000000000000000000000000000000000; // D (0x0000040800000000) 
//    12'h72d : LOC <=          63'b000000000000000000010000000100000000000000000000000000000000000; // D (0x0000080800000000) 
//    12'hd27 : LOC <=          63'b000000000000000000100000000100000000000000000000000000000000000; // D (0x0000100800000000) 
//    12'hc0a : LOC <=          63'b000000000000000001000000000100000000000000000000000000000000000; // D (0x0000200800000000) 
//    12'he50 : LOC <=          63'b000000000000000010000000000100000000000000000000000000000000000; // D (0x0000400800000000) 
//    12'hae4 : LOC <=          63'b000000000000000100000000000100000000000000000000000000000000000; // D (0x0000800800000000) 
//    12'h38c : LOC <=          63'b000000000000001000000000000100000000000000000000000000000000000; // D (0x0001000800000000) 
//    12'h465 : LOC <=          63'b000000000000010000000000000100000000000000000000000000000000000; // D (0x0002000800000000) 
//    12'hbb7 : LOC <=          63'b000000000000100000000000000100000000000000000000000000000000000; // D (0x0004000800000000) 
//    12'h12a : LOC <=          63'b000000000001000000000000000100000000000000000000000000000000000; // D (0x0008000800000000) 
//    12'h129 : LOC <=          63'b000000000010000000000000000100000000000000000000000000000000000; // D (0x0010000800000000) 
//    12'h12f : LOC <=          63'b000000000100000000000000000100000000000000000000000000000000000; // D (0x0020000800000000) 
//    12'h123 : LOC <=          63'b000000001000000000000000000100000000000000000000000000000000000; // D (0x0040000800000000) 
//    12'h13b : LOC <=          63'b000000010000000000000000000100000000000000000000000000000000000; // D (0x0080000800000000) 
//    12'h10b : LOC <=          63'b000000100000000000000000000100000000000000000000000000000000000; // D (0x0100000800000000) 
//    12'h16b : LOC <=          63'b000001000000000000000000000100000000000000000000000000000000000; // D (0x0200000800000000) 
//    12'h1ab : LOC <=          63'b000010000000000000000000000100000000000000000000000000000000000; // D (0x0400000800000000) 
//    12'h02b : LOC <=          63'b000100000000000000000000000100000000000000000000000000000000000; // D (0x0800000800000000) 
//    12'h32b : LOC <=          63'b001000000000000000000000000100000000000000000000000000000000000; // D (0x1000000800000000) 
//    12'h52b : LOC <=          63'b010000000000000000000000000100000000000000000000000000000000000; // D (0x2000000800000000) 
//    12'h92b : LOC <=          63'b100000000000000000000000000100000000000000000000000000000000000; // D (0x4000000800000000) 
    12'h76f : LOC <=          63'b000000000000000000000000001000000000000000000000000000000000001; // D (0x0000001000000001) 
    12'h824 : LOC <=          63'b000000000000000000000000001000000000000000000000000000000000010; // D (0x0000001000000002) 
    12'h38b : LOC <=          63'b000000000000000000000000001000000000000000000000000000000000100; // D (0x0000001000000004) 
    12'h1ec : LOC <=          63'b000000000000000000000000001000000000000000000000000000000001000; // D (0x0000001000000008) 
    12'h522 : LOC <=          63'b000000000000000000000000001000000000000000000000000000000010000; // D (0x0000001000000010) 
    12'hcbe : LOC <=          63'b000000000000000000000000001000000000000000000000000000000100000; // D (0x0000001000000020) 
    12'habf : LOC <=          63'b000000000000000000000000001000000000000000000000000000001000000; // D (0x0000001000000040) 
    12'h6bd : LOC <=          63'b000000000000000000000000001000000000000000000000000000010000000; // D (0x0000001000000080) 
    12'hb80 : LOC <=          63'b000000000000000000000000001000000000000000000000000000100000000; // D (0x0000001000000100) 
    12'h4c3 : LOC <=          63'b000000000000000000000000001000000000000000000000000001000000000; // D (0x0000001000000200) 
    12'hf7c : LOC <=          63'b000000000000000000000000001000000000000000000000000010000000000; // D (0x0000001000000400) 
    12'hd3b : LOC <=          63'b000000000000000000000000001000000000000000000000000100000000000; // D (0x0000001000000800) 
    12'h9b5 : LOC <=          63'b000000000000000000000000001000000000000000000000001000000000000; // D (0x0000001000001000) 
    12'h0a9 : LOC <=          63'b000000000000000000000000001000000000000000000000010000000000000; // D (0x0000001000002000) 
    12'h7a8 : LOC <=          63'b000000000000000000000000001000000000000000000000100000000000000; // D (0x0000001000004000) 
    12'h9aa : LOC <=          63'b000000000000000000000000001000000000000000000001000000000000000; // D (0x0000001000008000) 
    12'h097 : LOC <=          63'b000000000000000000000000001000000000000000000010000000000000000; // D (0x0000001000010000) 
    12'h7d4 : LOC <=          63'b000000000000000000000000001000000000000000000100000000000000000; // D (0x0000001000020000) 
    12'h952 : LOC <=          63'b000000000000000000000000001000000000000000001000000000000000000; // D (0x0000001000040000) 
    12'h167 : LOC <=          63'b000000000000000000000000001000000000000000010000000000000000000; // D (0x0000001000080000) 
    12'h434 : LOC <=          63'b000000000000000000000000001000000000000000100000000000000000000; // D (0x0000001000100000) 
    12'he92 : LOC <=          63'b000000000000000000000000001000000000000001000000000000000000000; // D (0x0000001000200000) 
    12'hee7 : LOC <=          63'b000000000000000000000000001000000000000010000000000000000000000; // D (0x0000001000400000) 
    12'he0d : LOC <=          63'b000000000000000000000000001000000000000100000000000000000000000; // D (0x0000001000800000) 
    12'hfd9 : LOC <=          63'b000000000000000000000000001000000000001000000000000000000000000; // D (0x0000001001000000) 
    12'hc71 : LOC <=          63'b000000000000000000000000001000000000010000000000000000000000000; // D (0x0000001002000000) 
    12'hb21 : LOC <=          63'b000000000000000000000000001000000000100000000000000000000000000; // D (0x0000001004000000) 
    12'h581 : LOC <=          63'b000000000000000000000000001000000001000000000000000000000000000; // D (0x0000001008000000) 
    12'hdf8 : LOC <=          63'b000000000000000000000000001000000010000000000000000000000000000; // D (0x0000001010000000) 
    12'h833 : LOC <=          63'b000000000000000000000000001000000100000000000000000000000000000; // D (0x0000001020000000) 
    12'h3a5 : LOC <=          63'b000000000000000000000000001000001000000000000000000000000000000; // D (0x0000001040000000) 
    12'h1b0 : LOC <=          63'b000000000000000000000000001000010000000000000000000000000000000; // D (0x0000001080000000) 
    12'h59a : LOC <=          63'b000000000000000000000000001000100000000000000000000000000000000; // D (0x0000001100000000) 
    12'hdce : LOC <=          63'b000000000000000000000000001001000000000000000000000000000000000; // D (0x0000001200000000) 
    12'h85f : LOC <=          63'b000000000000000000000000001010000000000000000000000000000000000; // D (0x0000001400000000) 
    12'h37d : LOC <=          63'b000000000000000000000000001100000000000000000000000000000000000; // D (0x0000001800000000) 
    12'h256 : LOC <=          63'b000000000000000000000000001000000000000000000000000000000000000; // S (0x0000001000000000) 
//    12'h6fa : LOC <=          63'b000000000000000000000000011000000000000000000000000000000000000; // D (0x0000003000000000) 
//    12'hb0e : LOC <=          63'b000000000000000000000000101000000000000000000000000000000000000; // D (0x0000005000000000) 
//    12'h5df : LOC <=          63'b000000000000000000000001001000000000000000000000000000000000000; // D (0x0000009000000000) 
//    12'hd44 : LOC <=          63'b000000000000000000000010001000000000000000000000000000000000000; // D (0x0000011000000000) 
//    12'h94b : LOC <=          63'b000000000000000000000100001000000000000000000000000000000000000; // D (0x0000021000000000) 
//    12'h155 : LOC <=          63'b000000000000000000001000001000000000000000000000000000000000000; // D (0x0000041000000000) 
//    12'h450 : LOC <=          63'b000000000000000000010000001000000000000000000000000000000000000; // D (0x0000081000000000) 
//    12'he5a : LOC <=          63'b000000000000000000100000001000000000000000000000000000000000000; // D (0x0000101000000000) 
//    12'hf77 : LOC <=          63'b000000000000000001000000001000000000000000000000000000000000000; // D (0x0000201000000000) 
//    12'hd2d : LOC <=          63'b000000000000000010000000001000000000000000000000000000000000000; // D (0x0000401000000000) 
//    12'h999 : LOC <=          63'b000000000000000100000000001000000000000000000000000000000000000; // D (0x0000801000000000) 
//    12'h0f1 : LOC <=          63'b000000000000001000000000001000000000000000000000000000000000000; // D (0x0001001000000000) 
//    12'h718 : LOC <=          63'b000000000000010000000000001000000000000000000000000000000000000; // D (0x0002001000000000) 
//    12'h8ca : LOC <=          63'b000000000000100000000000001000000000000000000000000000000000000; // D (0x0004001000000000) 
//    12'h257 : LOC <=          63'b000000000001000000000000001000000000000000000000000000000000000; // D (0x0008001000000000) 
//    12'h254 : LOC <=          63'b000000000010000000000000001000000000000000000000000000000000000; // D (0x0010001000000000) 
//    12'h252 : LOC <=          63'b000000000100000000000000001000000000000000000000000000000000000; // D (0x0020001000000000) 
//    12'h25e : LOC <=          63'b000000001000000000000000001000000000000000000000000000000000000; // D (0x0040001000000000) 
//    12'h246 : LOC <=          63'b000000010000000000000000001000000000000000000000000000000000000; // D (0x0080001000000000) 
//    12'h276 : LOC <=          63'b000000100000000000000000001000000000000000000000000000000000000; // D (0x0100001000000000) 
//    12'h216 : LOC <=          63'b000001000000000000000000001000000000000000000000000000000000000; // D (0x0200001000000000) 
//    12'h2d6 : LOC <=          63'b000010000000000000000000001000000000000000000000000000000000000; // D (0x0400001000000000) 
//    12'h356 : LOC <=          63'b000100000000000000000000001000000000000000000000000000000000000; // D (0x0800001000000000) 
//    12'h056 : LOC <=          63'b001000000000000000000000001000000000000000000000000000000000000; // D (0x1000001000000000) 
//    12'h656 : LOC <=          63'b010000000000000000000000001000000000000000000000000000000000000; // D (0x2000001000000000) 
//    12'ha56 : LOC <=          63'b100000000000000000000000001000000000000000000000000000000000000; // D (0x4000001000000000) 
    12'h195 : LOC <=          63'b000000000000000000000000010000000000000000000000000000000000001; // D (0x0000002000000001) 
    12'hede : LOC <=          63'b000000000000000000000000010000000000000000000000000000000000010; // D (0x0000002000000002) 
    12'h571 : LOC <=          63'b000000000000000000000000010000000000000000000000000000000000100; // D (0x0000002000000004) 
    12'h716 : LOC <=          63'b000000000000000000000000010000000000000000000000000000000001000; // D (0x0000002000000008) 
    12'h3d8 : LOC <=          63'b000000000000000000000000010000000000000000000000000000000010000; // D (0x0000002000000010) 
    12'ha44 : LOC <=          63'b000000000000000000000000010000000000000000000000000000000100000; // D (0x0000002000000020) 
    12'hc45 : LOC <=          63'b000000000000000000000000010000000000000000000000000000001000000; // D (0x0000002000000040) 
    12'h047 : LOC <=          63'b000000000000000000000000010000000000000000000000000000010000000; // D (0x0000002000000080) 
    12'hd7a : LOC <=          63'b000000000000000000000000010000000000000000000000000000100000000; // D (0x0000002000000100) 
    12'h239 : LOC <=          63'b000000000000000000000000010000000000000000000000000001000000000; // D (0x0000002000000200) 
    12'h986 : LOC <=          63'b000000000000000000000000010000000000000000000000000010000000000; // D (0x0000002000000400) 
    12'hbc1 : LOC <=          63'b000000000000000000000000010000000000000000000000000100000000000; // D (0x0000002000000800) 
    12'hf4f : LOC <=          63'b000000000000000000000000010000000000000000000000001000000000000; // D (0x0000002000001000) 
    12'h653 : LOC <=          63'b000000000000000000000000010000000000000000000000010000000000000; // D (0x0000002000002000) 
    12'h152 : LOC <=          63'b000000000000000000000000010000000000000000000000100000000000000; // D (0x0000002000004000) 
    12'hf50 : LOC <=          63'b000000000000000000000000010000000000000000000001000000000000000; // D (0x0000002000008000) 
    12'h66d : LOC <=          63'b000000000000000000000000010000000000000000000010000000000000000; // D (0x0000002000010000) 
    12'h12e : LOC <=          63'b000000000000000000000000010000000000000000000100000000000000000; // D (0x0000002000020000) 
    12'hfa8 : LOC <=          63'b000000000000000000000000010000000000000000001000000000000000000; // D (0x0000002000040000) 
    12'h79d : LOC <=          63'b000000000000000000000000010000000000000000010000000000000000000; // D (0x0000002000080000) 
    12'h2ce : LOC <=          63'b000000000000000000000000010000000000000000100000000000000000000; // D (0x0000002000100000) 
    12'h868 : LOC <=          63'b000000000000000000000000010000000000000001000000000000000000000; // D (0x0000002000200000) 
    12'h81d : LOC <=          63'b000000000000000000000000010000000000000010000000000000000000000; // D (0x0000002000400000) 
    12'h8f7 : LOC <=          63'b000000000000000000000000010000000000000100000000000000000000000; // D (0x0000002000800000) 
    12'h923 : LOC <=          63'b000000000000000000000000010000000000001000000000000000000000000; // D (0x0000002001000000) 
    12'ha8b : LOC <=          63'b000000000000000000000000010000000000010000000000000000000000000; // D (0x0000002002000000) 
    12'hddb : LOC <=          63'b000000000000000000000000010000000000100000000000000000000000000; // D (0x0000002004000000) 
    12'h37b : LOC <=          63'b000000000000000000000000010000000001000000000000000000000000000; // D (0x0000002008000000) 
    12'hb02 : LOC <=          63'b000000000000000000000000010000000010000000000000000000000000000; // D (0x0000002010000000) 
    12'hec9 : LOC <=          63'b000000000000000000000000010000000100000000000000000000000000000; // D (0x0000002020000000) 
    12'h55f : LOC <=          63'b000000000000000000000000010000001000000000000000000000000000000; // D (0x0000002040000000) 
    12'h74a : LOC <=          63'b000000000000000000000000010000010000000000000000000000000000000; // D (0x0000002080000000) 
    12'h360 : LOC <=          63'b000000000000000000000000010000100000000000000000000000000000000; // D (0x0000002100000000) 
    12'hb34 : LOC <=          63'b000000000000000000000000010001000000000000000000000000000000000; // D (0x0000002200000000) 
    12'hea5 : LOC <=          63'b000000000000000000000000010010000000000000000000000000000000000; // D (0x0000002400000000) 
    12'h587 : LOC <=          63'b000000000000000000000000010100000000000000000000000000000000000; // D (0x0000002800000000) 
    12'h6fa : LOC <=          63'b000000000000000000000000011000000000000000000000000000000000000; // D (0x0000003000000000) 
    12'h4ac : LOC <=          63'b000000000000000000000000010000000000000000000000000000000000000; // S (0x0000002000000000) 
//    12'hdf4 : LOC <=          63'b000000000000000000000000110000000000000000000000000000000000000; // D (0x0000006000000000) 
//    12'h325 : LOC <=          63'b000000000000000000000001010000000000000000000000000000000000000; // D (0x000000a000000000) 
//    12'hbbe : LOC <=          63'b000000000000000000000010010000000000000000000000000000000000000; // D (0x0000012000000000) 
//    12'hfb1 : LOC <=          63'b000000000000000000000100010000000000000000000000000000000000000; // D (0x0000022000000000) 
//    12'h7af : LOC <=          63'b000000000000000000001000010000000000000000000000000000000000000; // D (0x0000042000000000) 
//    12'h2aa : LOC <=          63'b000000000000000000010000010000000000000000000000000000000000000; // D (0x0000082000000000) 
//    12'h8a0 : LOC <=          63'b000000000000000000100000010000000000000000000000000000000000000; // D (0x0000102000000000) 
//    12'h98d : LOC <=          63'b000000000000000001000000010000000000000000000000000000000000000; // D (0x0000202000000000) 
//    12'hbd7 : LOC <=          63'b000000000000000010000000010000000000000000000000000000000000000; // D (0x0000402000000000) 
//    12'hf63 : LOC <=          63'b000000000000000100000000010000000000000000000000000000000000000; // D (0x0000802000000000) 
//    12'h60b : LOC <=          63'b000000000000001000000000010000000000000000000000000000000000000; // D (0x0001002000000000) 
//    12'h1e2 : LOC <=          63'b000000000000010000000000010000000000000000000000000000000000000; // D (0x0002002000000000) 
//    12'he30 : LOC <=          63'b000000000000100000000000010000000000000000000000000000000000000; // D (0x0004002000000000) 
//    12'h4ad : LOC <=          63'b000000000001000000000000010000000000000000000000000000000000000; // D (0x0008002000000000) 
//    12'h4ae : LOC <=          63'b000000000010000000000000010000000000000000000000000000000000000; // D (0x0010002000000000) 
//    12'h4a8 : LOC <=          63'b000000000100000000000000010000000000000000000000000000000000000; // D (0x0020002000000000) 
//    12'h4a4 : LOC <=          63'b000000001000000000000000010000000000000000000000000000000000000; // D (0x0040002000000000) 
//    12'h4bc : LOC <=          63'b000000010000000000000000010000000000000000000000000000000000000; // D (0x0080002000000000) 
//    12'h48c : LOC <=          63'b000000100000000000000000010000000000000000000000000000000000000; // D (0x0100002000000000) 
//    12'h4ec : LOC <=          63'b000001000000000000000000010000000000000000000000000000000000000; // D (0x0200002000000000) 
//    12'h42c : LOC <=          63'b000010000000000000000000010000000000000000000000000000000000000; // D (0x0400002000000000) 
//    12'h5ac : LOC <=          63'b000100000000000000000000010000000000000000000000000000000000000; // D (0x0800002000000000) 
//    12'h6ac : LOC <=          63'b001000000000000000000000010000000000000000000000000000000000000; // D (0x1000002000000000) 
//    12'h0ac : LOC <=          63'b010000000000000000000000010000000000000000000000000000000000000; // D (0x2000002000000000) 
//    12'hcac : LOC <=          63'b100000000000000000000000010000000000000000000000000000000000000; // D (0x4000002000000000) 
    12'hc61 : LOC <=          63'b000000000000000000000000100000000000000000000000000000000000001; // D (0x0000004000000001) 
    12'h32a : LOC <=          63'b000000000000000000000000100000000000000000000000000000000000010; // D (0x0000004000000002) 
    12'h885 : LOC <=          63'b000000000000000000000000100000000000000000000000000000000000100; // D (0x0000004000000004) 
    12'hae2 : LOC <=          63'b000000000000000000000000100000000000000000000000000000000001000; // D (0x0000004000000008) 
    12'he2c : LOC <=          63'b000000000000000000000000100000000000000000000000000000000010000; // D (0x0000004000000010) 
    12'h7b0 : LOC <=          63'b000000000000000000000000100000000000000000000000000000000100000; // D (0x0000004000000020) 
    12'h1b1 : LOC <=          63'b000000000000000000000000100000000000000000000000000000001000000; // D (0x0000004000000040) 
    12'hdb3 : LOC <=          63'b000000000000000000000000100000000000000000000000000000010000000; // D (0x0000004000000080) 
    12'h08e : LOC <=          63'b000000000000000000000000100000000000000000000000000000100000000; // D (0x0000004000000100) 
    12'hfcd : LOC <=          63'b000000000000000000000000100000000000000000000000000001000000000; // D (0x0000004000000200) 
    12'h472 : LOC <=          63'b000000000000000000000000100000000000000000000000000010000000000; // D (0x0000004000000400) 
    12'h635 : LOC <=          63'b000000000000000000000000100000000000000000000000000100000000000; // D (0x0000004000000800) 
    12'h2bb : LOC <=          63'b000000000000000000000000100000000000000000000000001000000000000; // D (0x0000004000001000) 
    12'hba7 : LOC <=          63'b000000000000000000000000100000000000000000000000010000000000000; // D (0x0000004000002000) 
    12'hca6 : LOC <=          63'b000000000000000000000000100000000000000000000000100000000000000; // D (0x0000004000004000) 
    12'h2a4 : LOC <=          63'b000000000000000000000000100000000000000000000001000000000000000; // D (0x0000004000008000) 
    12'hb99 : LOC <=          63'b000000000000000000000000100000000000000000000010000000000000000; // D (0x0000004000010000) 
    12'hcda : LOC <=          63'b000000000000000000000000100000000000000000000100000000000000000; // D (0x0000004000020000) 
    12'h25c : LOC <=          63'b000000000000000000000000100000000000000000001000000000000000000; // D (0x0000004000040000) 
    12'ha69 : LOC <=          63'b000000000000000000000000100000000000000000010000000000000000000; // D (0x0000004000080000) 
    12'hf3a : LOC <=          63'b000000000000000000000000100000000000000000100000000000000000000; // D (0x0000004000100000) 
    12'h59c : LOC <=          63'b000000000000000000000000100000000000000001000000000000000000000; // D (0x0000004000200000) 
    12'h5e9 : LOC <=          63'b000000000000000000000000100000000000000010000000000000000000000; // D (0x0000004000400000) 
    12'h503 : LOC <=          63'b000000000000000000000000100000000000000100000000000000000000000; // D (0x0000004000800000) 
    12'h4d7 : LOC <=          63'b000000000000000000000000100000000000001000000000000000000000000; // D (0x0000004001000000) 
    12'h77f : LOC <=          63'b000000000000000000000000100000000000010000000000000000000000000; // D (0x0000004002000000) 
    12'h02f : LOC <=          63'b000000000000000000000000100000000000100000000000000000000000000; // D (0x0000004004000000) 
    12'he8f : LOC <=          63'b000000000000000000000000100000000001000000000000000000000000000; // D (0x0000004008000000) 
    12'h6f6 : LOC <=          63'b000000000000000000000000100000000010000000000000000000000000000; // D (0x0000004010000000) 
    12'h33d : LOC <=          63'b000000000000000000000000100000000100000000000000000000000000000; // D (0x0000004020000000) 
    12'h8ab : LOC <=          63'b000000000000000000000000100000001000000000000000000000000000000; // D (0x0000004040000000) 
    12'habe : LOC <=          63'b000000000000000000000000100000010000000000000000000000000000000; // D (0x0000004080000000) 
    12'he94 : LOC <=          63'b000000000000000000000000100000100000000000000000000000000000000; // D (0x0000004100000000) 
    12'h6c0 : LOC <=          63'b000000000000000000000000100001000000000000000000000000000000000; // D (0x0000004200000000) 
    12'h351 : LOC <=          63'b000000000000000000000000100010000000000000000000000000000000000; // D (0x0000004400000000) 
    12'h873 : LOC <=          63'b000000000000000000000000100100000000000000000000000000000000000; // D (0x0000004800000000) 
    12'hb0e : LOC <=          63'b000000000000000000000000101000000000000000000000000000000000000; // D (0x0000005000000000) 
    12'hdf4 : LOC <=          63'b000000000000000000000000110000000000000000000000000000000000000; // D (0x0000006000000000) 
    12'h958 : LOC <=          63'b000000000000000000000000100000000000000000000000000000000000000; // S (0x0000004000000000) 
//    12'hed1 : LOC <=          63'b000000000000000000000001100000000000000000000000000000000000000; // D (0x000000c000000000) 
//    12'h64a : LOC <=          63'b000000000000000000000010100000000000000000000000000000000000000; // D (0x0000014000000000) 
//    12'h245 : LOC <=          63'b000000000000000000000100100000000000000000000000000000000000000; // D (0x0000024000000000) 
//    12'ha5b : LOC <=          63'b000000000000000000001000100000000000000000000000000000000000000; // D (0x0000044000000000) 
//    12'hf5e : LOC <=          63'b000000000000000000010000100000000000000000000000000000000000000; // D (0x0000084000000000) 
//    12'h554 : LOC <=          63'b000000000000000000100000100000000000000000000000000000000000000; // D (0x0000104000000000) 
//    12'h479 : LOC <=          63'b000000000000000001000000100000000000000000000000000000000000000; // D (0x0000204000000000) 
//    12'h623 : LOC <=          63'b000000000000000010000000100000000000000000000000000000000000000; // D (0x0000404000000000) 
//    12'h297 : LOC <=          63'b000000000000000100000000100000000000000000000000000000000000000; // D (0x0000804000000000) 
//    12'hbff : LOC <=          63'b000000000000001000000000100000000000000000000000000000000000000; // D (0x0001004000000000) 
//    12'hc16 : LOC <=          63'b000000000000010000000000100000000000000000000000000000000000000; // D (0x0002004000000000) 
//    12'h3c4 : LOC <=          63'b000000000000100000000000100000000000000000000000000000000000000; // D (0x0004004000000000) 
//    12'h959 : LOC <=          63'b000000000001000000000000100000000000000000000000000000000000000; // D (0x0008004000000000) 
//    12'h95a : LOC <=          63'b000000000010000000000000100000000000000000000000000000000000000; // D (0x0010004000000000) 
//    12'h95c : LOC <=          63'b000000000100000000000000100000000000000000000000000000000000000; // D (0x0020004000000000) 
//    12'h950 : LOC <=          63'b000000001000000000000000100000000000000000000000000000000000000; // D (0x0040004000000000) 
//    12'h948 : LOC <=          63'b000000010000000000000000100000000000000000000000000000000000000; // D (0x0080004000000000) 
//    12'h978 : LOC <=          63'b000000100000000000000000100000000000000000000000000000000000000; // D (0x0100004000000000) 
//    12'h918 : LOC <=          63'b000001000000000000000000100000000000000000000000000000000000000; // D (0x0200004000000000) 
//    12'h9d8 : LOC <=          63'b000010000000000000000000100000000000000000000000000000000000000; // D (0x0400004000000000) 
//    12'h858 : LOC <=          63'b000100000000000000000000100000000000000000000000000000000000000; // D (0x0800004000000000) 
//    12'hb58 : LOC <=          63'b001000000000000000000000100000000000000000000000000000000000000; // D (0x1000004000000000) 
//    12'hd58 : LOC <=          63'b010000000000000000000000100000000000000000000000000000000000000; // D (0x2000004000000000) 
//    12'h158 : LOC <=          63'b100000000000000000000000100000000000000000000000000000000000000; // D (0x4000004000000000) 
    12'h2b0 : LOC <=          63'b000000000000000000000001000000000000000000000000000000000000001; // D (0x0000008000000001) 
    12'hdfb : LOC <=          63'b000000000000000000000001000000000000000000000000000000000000010; // D (0x0000008000000002) 
    12'h654 : LOC <=          63'b000000000000000000000001000000000000000000000000000000000000100; // D (0x0000008000000004) 
    12'h433 : LOC <=          63'b000000000000000000000001000000000000000000000000000000000001000; // D (0x0000008000000008) 
    12'h0fd : LOC <=          63'b000000000000000000000001000000000000000000000000000000000010000; // D (0x0000008000000010) 
    12'h961 : LOC <=          63'b000000000000000000000001000000000000000000000000000000000100000; // D (0x0000008000000020) 
    12'hf60 : LOC <=          63'b000000000000000000000001000000000000000000000000000000001000000; // D (0x0000008000000040) 
    12'h362 : LOC <=          63'b000000000000000000000001000000000000000000000000000000010000000; // D (0x0000008000000080) 
    12'he5f : LOC <=          63'b000000000000000000000001000000000000000000000000000000100000000; // D (0x0000008000000100) 
    12'h11c : LOC <=          63'b000000000000000000000001000000000000000000000000000001000000000; // D (0x0000008000000200) 
    12'haa3 : LOC <=          63'b000000000000000000000001000000000000000000000000000010000000000; // D (0x0000008000000400) 
    12'h8e4 : LOC <=          63'b000000000000000000000001000000000000000000000000000100000000000; // D (0x0000008000000800) 
    12'hc6a : LOC <=          63'b000000000000000000000001000000000000000000000000001000000000000; // D (0x0000008000001000) 
    12'h576 : LOC <=          63'b000000000000000000000001000000000000000000000000010000000000000; // D (0x0000008000002000) 
    12'h277 : LOC <=          63'b000000000000000000000001000000000000000000000000100000000000000; // D (0x0000008000004000) 
    12'hc75 : LOC <=          63'b000000000000000000000001000000000000000000000001000000000000000; // D (0x0000008000008000) 
    12'h548 : LOC <=          63'b000000000000000000000001000000000000000000000010000000000000000; // D (0x0000008000010000) 
    12'h20b : LOC <=          63'b000000000000000000000001000000000000000000000100000000000000000; // D (0x0000008000020000) 
    12'hc8d : LOC <=          63'b000000000000000000000001000000000000000000001000000000000000000; // D (0x0000008000040000) 
    12'h4b8 : LOC <=          63'b000000000000000000000001000000000000000000010000000000000000000; // D (0x0000008000080000) 
    12'h1eb : LOC <=          63'b000000000000000000000001000000000000000000100000000000000000000; // D (0x0000008000100000) 
    12'hb4d : LOC <=          63'b000000000000000000000001000000000000000001000000000000000000000; // D (0x0000008000200000) 
    12'hb38 : LOC <=          63'b000000000000000000000001000000000000000010000000000000000000000; // D (0x0000008000400000) 
    12'hbd2 : LOC <=          63'b000000000000000000000001000000000000000100000000000000000000000; // D (0x0000008000800000) 
    12'ha06 : LOC <=          63'b000000000000000000000001000000000000001000000000000000000000000; // D (0x0000008001000000) 
    12'h9ae : LOC <=          63'b000000000000000000000001000000000000010000000000000000000000000; // D (0x0000008002000000) 
    12'hefe : LOC <=          63'b000000000000000000000001000000000000100000000000000000000000000; // D (0x0000008004000000) 
    12'h05e : LOC <=          63'b000000000000000000000001000000000001000000000000000000000000000; // D (0x0000008008000000) 
    12'h827 : LOC <=          63'b000000000000000000000001000000000010000000000000000000000000000; // D (0x0000008010000000) 
    12'hdec : LOC <=          63'b000000000000000000000001000000000100000000000000000000000000000; // D (0x0000008020000000) 
    12'h67a : LOC <=          63'b000000000000000000000001000000001000000000000000000000000000000; // D (0x0000008040000000) 
    12'h46f : LOC <=          63'b000000000000000000000001000000010000000000000000000000000000000; // D (0x0000008080000000) 
    12'h045 : LOC <=          63'b000000000000000000000001000000100000000000000000000000000000000; // D (0x0000008100000000) 
    12'h811 : LOC <=          63'b000000000000000000000001000001000000000000000000000000000000000; // D (0x0000008200000000) 
    12'hd80 : LOC <=          63'b000000000000000000000001000010000000000000000000000000000000000; // D (0x0000008400000000) 
    12'h6a2 : LOC <=          63'b000000000000000000000001000100000000000000000000000000000000000; // D (0x0000008800000000) 
    12'h5df : LOC <=          63'b000000000000000000000001001000000000000000000000000000000000000; // D (0x0000009000000000) 
    12'h325 : LOC <=          63'b000000000000000000000001010000000000000000000000000000000000000; // D (0x000000a000000000) 
    12'hed1 : LOC <=          63'b000000000000000000000001100000000000000000000000000000000000000; // D (0x000000c000000000) 
    12'h789 : LOC <=          63'b000000000000000000000001000000000000000000000000000000000000000; // S (0x0000008000000000) 
//    12'h89b : LOC <=          63'b000000000000000000000011000000000000000000000000000000000000000; // D (0x0000018000000000) 
//    12'hc94 : LOC <=          63'b000000000000000000000101000000000000000000000000000000000000000; // D (0x0000028000000000) 
//    12'h48a : LOC <=          63'b000000000000000000001001000000000000000000000000000000000000000; // D (0x0000048000000000) 
//    12'h18f : LOC <=          63'b000000000000000000010001000000000000000000000000000000000000000; // D (0x0000088000000000) 
//    12'hb85 : LOC <=          63'b000000000000000000100001000000000000000000000000000000000000000; // D (0x0000108000000000) 
//    12'haa8 : LOC <=          63'b000000000000000001000001000000000000000000000000000000000000000; // D (0x0000208000000000) 
//    12'h8f2 : LOC <=          63'b000000000000000010000001000000000000000000000000000000000000000; // D (0x0000408000000000) 
//    12'hc46 : LOC <=          63'b000000000000000100000001000000000000000000000000000000000000000; // D (0x0000808000000000) 
//    12'h52e : LOC <=          63'b000000000000001000000001000000000000000000000000000000000000000; // D (0x0001008000000000) 
//    12'h2c7 : LOC <=          63'b000000000000010000000001000000000000000000000000000000000000000; // D (0x0002008000000000) 
//    12'hd15 : LOC <=          63'b000000000000100000000001000000000000000000000000000000000000000; // D (0x0004008000000000) 
//    12'h788 : LOC <=          63'b000000000001000000000001000000000000000000000000000000000000000; // D (0x0008008000000000) 
//    12'h78b : LOC <=          63'b000000000010000000000001000000000000000000000000000000000000000; // D (0x0010008000000000) 
//    12'h78d : LOC <=          63'b000000000100000000000001000000000000000000000000000000000000000; // D (0x0020008000000000) 
//    12'h781 : LOC <=          63'b000000001000000000000001000000000000000000000000000000000000000; // D (0x0040008000000000) 
//    12'h799 : LOC <=          63'b000000010000000000000001000000000000000000000000000000000000000; // D (0x0080008000000000) 
//    12'h7a9 : LOC <=          63'b000000100000000000000001000000000000000000000000000000000000000; // D (0x0100008000000000) 
//    12'h7c9 : LOC <=          63'b000001000000000000000001000000000000000000000000000000000000000; // D (0x0200008000000000) 
//    12'h709 : LOC <=          63'b000010000000000000000001000000000000000000000000000000000000000; // D (0x0400008000000000) 
//    12'h689 : LOC <=          63'b000100000000000000000001000000000000000000000000000000000000000; // D (0x0800008000000000) 
//    12'h589 : LOC <=          63'b001000000000000000000001000000000000000000000000000000000000000; // D (0x1000008000000000) 
//    12'h389 : LOC <=          63'b010000000000000000000001000000000000000000000000000000000000000; // D (0x2000008000000000) 
//    12'hf89 : LOC <=          63'b100000000000000000000001000000000000000000000000000000000000000; // D (0x4000008000000000) 
    12'ha2b : LOC <=          63'b000000000000000000000010000000000000000000000000000000000000001; // D (0x0000010000000001) 
    12'h560 : LOC <=          63'b000000000000000000000010000000000000000000000000000000000000010; // D (0x0000010000000002) 
    12'hecf : LOC <=          63'b000000000000000000000010000000000000000000000000000000000000100; // D (0x0000010000000004) 
    12'hca8 : LOC <=          63'b000000000000000000000010000000000000000000000000000000000001000; // D (0x0000010000000008) 
    12'h866 : LOC <=          63'b000000000000000000000010000000000000000000000000000000000010000; // D (0x0000010000000010) 
    12'h1fa : LOC <=          63'b000000000000000000000010000000000000000000000000000000000100000; // D (0x0000010000000020) 
    12'h7fb : LOC <=          63'b000000000000000000000010000000000000000000000000000000001000000; // D (0x0000010000000040) 
    12'hbf9 : LOC <=          63'b000000000000000000000010000000000000000000000000000000010000000; // D (0x0000010000000080) 
    12'h6c4 : LOC <=          63'b000000000000000000000010000000000000000000000000000000100000000; // D (0x0000010000000100) 
    12'h987 : LOC <=          63'b000000000000000000000010000000000000000000000000000001000000000; // D (0x0000010000000200) 
    12'h238 : LOC <=          63'b000000000000000000000010000000000000000000000000000010000000000; // D (0x0000010000000400) 
    12'h07f : LOC <=          63'b000000000000000000000010000000000000000000000000000100000000000; // D (0x0000010000000800) 
    12'h4f1 : LOC <=          63'b000000000000000000000010000000000000000000000000001000000000000; // D (0x0000010000001000) 
    12'hded : LOC <=          63'b000000000000000000000010000000000000000000000000010000000000000; // D (0x0000010000002000) 
    12'haec : LOC <=          63'b000000000000000000000010000000000000000000000000100000000000000; // D (0x0000010000004000) 
    12'h4ee : LOC <=          63'b000000000000000000000010000000000000000000000001000000000000000; // D (0x0000010000008000) 
    12'hdd3 : LOC <=          63'b000000000000000000000010000000000000000000000010000000000000000; // D (0x0000010000010000) 
    12'ha90 : LOC <=          63'b000000000000000000000010000000000000000000000100000000000000000; // D (0x0000010000020000) 
    12'h416 : LOC <=          63'b000000000000000000000010000000000000000000001000000000000000000; // D (0x0000010000040000) 
    12'hc23 : LOC <=          63'b000000000000000000000010000000000000000000010000000000000000000; // D (0x0000010000080000) 
    12'h970 : LOC <=          63'b000000000000000000000010000000000000000000100000000000000000000; // D (0x0000010000100000) 
    12'h3d6 : LOC <=          63'b000000000000000000000010000000000000000001000000000000000000000; // D (0x0000010000200000) 
    12'h3a3 : LOC <=          63'b000000000000000000000010000000000000000010000000000000000000000; // D (0x0000010000400000) 
    12'h349 : LOC <=          63'b000000000000000000000010000000000000000100000000000000000000000; // D (0x0000010000800000) 
    12'h29d : LOC <=          63'b000000000000000000000010000000000000001000000000000000000000000; // D (0x0000010001000000) 
    12'h135 : LOC <=          63'b000000000000000000000010000000000000010000000000000000000000000; // D (0x0000010002000000) 
    12'h665 : LOC <=          63'b000000000000000000000010000000000000100000000000000000000000000; // D (0x0000010004000000) 
    12'h8c5 : LOC <=          63'b000000000000000000000010000000000001000000000000000000000000000; // D (0x0000010008000000) 
    12'h0bc : LOC <=          63'b000000000000000000000010000000000010000000000000000000000000000; // D (0x0000010010000000) 
    12'h577 : LOC <=          63'b000000000000000000000010000000000100000000000000000000000000000; // D (0x0000010020000000) 
    12'hee1 : LOC <=          63'b000000000000000000000010000000001000000000000000000000000000000; // D (0x0000010040000000) 
    12'hcf4 : LOC <=          63'b000000000000000000000010000000010000000000000000000000000000000; // D (0x0000010080000000) 
    12'h8de : LOC <=          63'b000000000000000000000010000000100000000000000000000000000000000; // D (0x0000010100000000) 
    12'h08a : LOC <=          63'b000000000000000000000010000001000000000000000000000000000000000; // D (0x0000010200000000) 
    12'h51b : LOC <=          63'b000000000000000000000010000010000000000000000000000000000000000; // D (0x0000010400000000) 
    12'he39 : LOC <=          63'b000000000000000000000010000100000000000000000000000000000000000; // D (0x0000010800000000) 
    12'hd44 : LOC <=          63'b000000000000000000000010001000000000000000000000000000000000000; // D (0x0000011000000000) 
    12'hbbe : LOC <=          63'b000000000000000000000010010000000000000000000000000000000000000; // D (0x0000012000000000) 
    12'h64a : LOC <=          63'b000000000000000000000010100000000000000000000000000000000000000; // D (0x0000014000000000) 
    12'h89b : LOC <=          63'b000000000000000000000011000000000000000000000000000000000000000; // D (0x0000018000000000) 
    12'hf12 : LOC <=          63'b000000000000000000000010000000000000000000000000000000000000000; // S (0x0000010000000000) 
//    12'h40f : LOC <=          63'b000000000000000000000110000000000000000000000000000000000000000; // D (0x0000030000000000) 
//    12'hc11 : LOC <=          63'b000000000000000000001010000000000000000000000000000000000000000; // D (0x0000050000000000) 
//    12'h914 : LOC <=          63'b000000000000000000010010000000000000000000000000000000000000000; // D (0x0000090000000000) 
//    12'h31e : LOC <=          63'b000000000000000000100010000000000000000000000000000000000000000; // D (0x0000110000000000) 
//    12'h233 : LOC <=          63'b000000000000000001000010000000000000000000000000000000000000000; // D (0x0000210000000000) 
//    12'h069 : LOC <=          63'b000000000000000010000010000000000000000000000000000000000000000; // D (0x0000410000000000) 
//    12'h4dd : LOC <=          63'b000000000000000100000010000000000000000000000000000000000000000; // D (0x0000810000000000) 
//    12'hdb5 : LOC <=          63'b000000000000001000000010000000000000000000000000000000000000000; // D (0x0001010000000000) 
//    12'ha5c : LOC <=          63'b000000000000010000000010000000000000000000000000000000000000000; // D (0x0002010000000000) 
//    12'h58e : LOC <=          63'b000000000000100000000010000000000000000000000000000000000000000; // D (0x0004010000000000) 
//    12'hf13 : LOC <=          63'b000000000001000000000010000000000000000000000000000000000000000; // D (0x0008010000000000) 
//    12'hf10 : LOC <=          63'b000000000010000000000010000000000000000000000000000000000000000; // D (0x0010010000000000) 
//    12'hf16 : LOC <=          63'b000000000100000000000010000000000000000000000000000000000000000; // D (0x0020010000000000) 
//    12'hf1a : LOC <=          63'b000000001000000000000010000000000000000000000000000000000000000; // D (0x0040010000000000) 
//    12'hf02 : LOC <=          63'b000000010000000000000010000000000000000000000000000000000000000; // D (0x0080010000000000) 
//    12'hf32 : LOC <=          63'b000000100000000000000010000000000000000000000000000000000000000; // D (0x0100010000000000) 
//    12'hf52 : LOC <=          63'b000001000000000000000010000000000000000000000000000000000000000; // D (0x0200010000000000) 
//    12'hf92 : LOC <=          63'b000010000000000000000010000000000000000000000000000000000000000; // D (0x0400010000000000) 
//    12'he12 : LOC <=          63'b000100000000000000000010000000000000000000000000000000000000000; // D (0x0800010000000000) 
//    12'hd12 : LOC <=          63'b001000000000000000000010000000000000000000000000000000000000000; // D (0x1000010000000000) 
//    12'hb12 : LOC <=          63'b010000000000000000000010000000000000000000000000000000000000000; // D (0x2000010000000000) 
//    12'h712 : LOC <=          63'b100000000000000000000010000000000000000000000000000000000000000; // D (0x4000010000000000) 
    12'he24 : LOC <=          63'b000000000000000000000100000000000000000000000000000000000000001; // D (0x0000020000000001) 
    12'h16f : LOC <=          63'b000000000000000000000100000000000000000000000000000000000000010; // D (0x0000020000000002) 
    12'hac0 : LOC <=          63'b000000000000000000000100000000000000000000000000000000000000100; // D (0x0000020000000004) 
    12'h8a7 : LOC <=          63'b000000000000000000000100000000000000000000000000000000000001000; // D (0x0000020000000008) 
    12'hc69 : LOC <=          63'b000000000000000000000100000000000000000000000000000000000010000; // D (0x0000020000000010) 
    12'h5f5 : LOC <=          63'b000000000000000000000100000000000000000000000000000000000100000; // D (0x0000020000000020) 
    12'h3f4 : LOC <=          63'b000000000000000000000100000000000000000000000000000000001000000; // D (0x0000020000000040) 
    12'hff6 : LOC <=          63'b000000000000000000000100000000000000000000000000000000010000000; // D (0x0000020000000080) 
    12'h2cb : LOC <=          63'b000000000000000000000100000000000000000000000000000000100000000; // D (0x0000020000000100) 
    12'hd88 : LOC <=          63'b000000000000000000000100000000000000000000000000000001000000000; // D (0x0000020000000200) 
    12'h637 : LOC <=          63'b000000000000000000000100000000000000000000000000000010000000000; // D (0x0000020000000400) 
    12'h470 : LOC <=          63'b000000000000000000000100000000000000000000000000000100000000000; // D (0x0000020000000800) 
    12'h0fe : LOC <=          63'b000000000000000000000100000000000000000000000000001000000000000; // D (0x0000020000001000) 
    12'h9e2 : LOC <=          63'b000000000000000000000100000000000000000000000000010000000000000; // D (0x0000020000002000) 
    12'hee3 : LOC <=          63'b000000000000000000000100000000000000000000000000100000000000000; // D (0x0000020000004000) 
    12'h0e1 : LOC <=          63'b000000000000000000000100000000000000000000000001000000000000000; // D (0x0000020000008000) 
    12'h9dc : LOC <=          63'b000000000000000000000100000000000000000000000010000000000000000; // D (0x0000020000010000) 
    12'he9f : LOC <=          63'b000000000000000000000100000000000000000000000100000000000000000; // D (0x0000020000020000) 
    12'h019 : LOC <=          63'b000000000000000000000100000000000000000000001000000000000000000; // D (0x0000020000040000) 
    12'h82c : LOC <=          63'b000000000000000000000100000000000000000000010000000000000000000; // D (0x0000020000080000) 
    12'hd7f : LOC <=          63'b000000000000000000000100000000000000000000100000000000000000000; // D (0x0000020000100000) 
    12'h7d9 : LOC <=          63'b000000000000000000000100000000000000000001000000000000000000000; // D (0x0000020000200000) 
    12'h7ac : LOC <=          63'b000000000000000000000100000000000000000010000000000000000000000; // D (0x0000020000400000) 
    12'h746 : LOC <=          63'b000000000000000000000100000000000000000100000000000000000000000; // D (0x0000020000800000) 
    12'h692 : LOC <=          63'b000000000000000000000100000000000000001000000000000000000000000; // D (0x0000020001000000) 
    12'h53a : LOC <=          63'b000000000000000000000100000000000000010000000000000000000000000; // D (0x0000020002000000) 
    12'h26a : LOC <=          63'b000000000000000000000100000000000000100000000000000000000000000; // D (0x0000020004000000) 
    12'hcca : LOC <=          63'b000000000000000000000100000000000001000000000000000000000000000; // D (0x0000020008000000) 
    12'h4b3 : LOC <=          63'b000000000000000000000100000000000010000000000000000000000000000; // D (0x0000020010000000) 
    12'h178 : LOC <=          63'b000000000000000000000100000000000100000000000000000000000000000; // D (0x0000020020000000) 
    12'haee : LOC <=          63'b000000000000000000000100000000001000000000000000000000000000000; // D (0x0000020040000000) 
    12'h8fb : LOC <=          63'b000000000000000000000100000000010000000000000000000000000000000; // D (0x0000020080000000) 
    12'hcd1 : LOC <=          63'b000000000000000000000100000000100000000000000000000000000000000; // D (0x0000020100000000) 
    12'h485 : LOC <=          63'b000000000000000000000100000001000000000000000000000000000000000; // D (0x0000020200000000) 
    12'h114 : LOC <=          63'b000000000000000000000100000010000000000000000000000000000000000; // D (0x0000020400000000) 
    12'ha36 : LOC <=          63'b000000000000000000000100000100000000000000000000000000000000000; // D (0x0000020800000000) 
    12'h94b : LOC <=          63'b000000000000000000000100001000000000000000000000000000000000000; // D (0x0000021000000000) 
    12'hfb1 : LOC <=          63'b000000000000000000000100010000000000000000000000000000000000000; // D (0x0000022000000000) 
    12'h245 : LOC <=          63'b000000000000000000000100100000000000000000000000000000000000000; // D (0x0000024000000000) 
    12'hc94 : LOC <=          63'b000000000000000000000101000000000000000000000000000000000000000; // D (0x0000028000000000) 
    12'h40f : LOC <=          63'b000000000000000000000110000000000000000000000000000000000000000; // D (0x0000030000000000) 
    12'hb1d : LOC <=          63'b000000000000000000000100000000000000000000000000000000000000000; // S (0x0000020000000000) 
//    12'h81e : LOC <=          63'b000000000000000000001100000000000000000000000000000000000000000; // D (0x0000060000000000) 
//    12'hd1b : LOC <=          63'b000000000000000000010100000000000000000000000000000000000000000; // D (0x00000a0000000000) 
//    12'h711 : LOC <=          63'b000000000000000000100100000000000000000000000000000000000000000; // D (0x0000120000000000) 
//    12'h63c : LOC <=          63'b000000000000000001000100000000000000000000000000000000000000000; // D (0x0000220000000000) 
//    12'h466 : LOC <=          63'b000000000000000010000100000000000000000000000000000000000000000; // D (0x0000420000000000) 
//    12'h0d2 : LOC <=          63'b000000000000000100000100000000000000000000000000000000000000000; // D (0x0000820000000000) 
//    12'h9ba : LOC <=          63'b000000000000001000000100000000000000000000000000000000000000000; // D (0x0001020000000000) 
//    12'he53 : LOC <=          63'b000000000000010000000100000000000000000000000000000000000000000; // D (0x0002020000000000) 
//    12'h181 : LOC <=          63'b000000000000100000000100000000000000000000000000000000000000000; // D (0x0004020000000000) 
//    12'hb1c : LOC <=          63'b000000000001000000000100000000000000000000000000000000000000000; // D (0x0008020000000000) 
//    12'hb1f : LOC <=          63'b000000000010000000000100000000000000000000000000000000000000000; // D (0x0010020000000000) 
//    12'hb19 : LOC <=          63'b000000000100000000000100000000000000000000000000000000000000000; // D (0x0020020000000000) 
//    12'hb15 : LOC <=          63'b000000001000000000000100000000000000000000000000000000000000000; // D (0x0040020000000000) 
//    12'hb0d : LOC <=          63'b000000010000000000000100000000000000000000000000000000000000000; // D (0x0080020000000000) 
//    12'hb3d : LOC <=          63'b000000100000000000000100000000000000000000000000000000000000000; // D (0x0100020000000000) 
//    12'hb5d : LOC <=          63'b000001000000000000000100000000000000000000000000000000000000000; // D (0x0200020000000000) 
//    12'hb9d : LOC <=          63'b000010000000000000000100000000000000000000000000000000000000000; // D (0x0400020000000000) 
//    12'ha1d : LOC <=          63'b000100000000000000000100000000000000000000000000000000000000000; // D (0x0800020000000000) 
//    12'h91d : LOC <=          63'b001000000000000000000100000000000000000000000000000000000000000; // D (0x1000020000000000) 
//    12'hf1d : LOC <=          63'b010000000000000000000100000000000000000000000000000000000000000; // D (0x2000020000000000) 
//    12'h31d : LOC <=          63'b100000000000000000000100000000000000000000000000000000000000000; // D (0x4000020000000000) 
    12'h63a : LOC <=          63'b000000000000000000001000000000000000000000000000000000000000001; // D (0x0000040000000001) 
    12'h971 : LOC <=          63'b000000000000000000001000000000000000000000000000000000000000010; // D (0x0000040000000002) 
    12'h2de : LOC <=          63'b000000000000000000001000000000000000000000000000000000000000100; // D (0x0000040000000004) 
    12'h0b9 : LOC <=          63'b000000000000000000001000000000000000000000000000000000000001000; // D (0x0000040000000008) 
    12'h477 : LOC <=          63'b000000000000000000001000000000000000000000000000000000000010000; // D (0x0000040000000010) 
    12'hdeb : LOC <=          63'b000000000000000000001000000000000000000000000000000000000100000; // D (0x0000040000000020) 
    12'hbea : LOC <=          63'b000000000000000000001000000000000000000000000000000000001000000; // D (0x0000040000000040) 
    12'h7e8 : LOC <=          63'b000000000000000000001000000000000000000000000000000000010000000; // D (0x0000040000000080) 
    12'had5 : LOC <=          63'b000000000000000000001000000000000000000000000000000000100000000; // D (0x0000040000000100) 
    12'h596 : LOC <=          63'b000000000000000000001000000000000000000000000000000001000000000; // D (0x0000040000000200) 
    12'he29 : LOC <=          63'b000000000000000000001000000000000000000000000000000010000000000; // D (0x0000040000000400) 
    12'hc6e : LOC <=          63'b000000000000000000001000000000000000000000000000000100000000000; // D (0x0000040000000800) 
    12'h8e0 : LOC <=          63'b000000000000000000001000000000000000000000000000001000000000000; // D (0x0000040000001000) 
    12'h1fc : LOC <=          63'b000000000000000000001000000000000000000000000000010000000000000; // D (0x0000040000002000) 
    12'h6fd : LOC <=          63'b000000000000000000001000000000000000000000000000100000000000000; // D (0x0000040000004000) 
    12'h8ff : LOC <=          63'b000000000000000000001000000000000000000000000001000000000000000; // D (0x0000040000008000) 
    12'h1c2 : LOC <=          63'b000000000000000000001000000000000000000000000010000000000000000; // D (0x0000040000010000) 
    12'h681 : LOC <=          63'b000000000000000000001000000000000000000000000100000000000000000; // D (0x0000040000020000) 
    12'h807 : LOC <=          63'b000000000000000000001000000000000000000000001000000000000000000; // D (0x0000040000040000) 
    12'h032 : LOC <=          63'b000000000000000000001000000000000000000000010000000000000000000; // D (0x0000040000080000) 
    12'h561 : LOC <=          63'b000000000000000000001000000000000000000000100000000000000000000; // D (0x0000040000100000) 
    12'hfc7 : LOC <=          63'b000000000000000000001000000000000000000001000000000000000000000; // D (0x0000040000200000) 
    12'hfb2 : LOC <=          63'b000000000000000000001000000000000000000010000000000000000000000; // D (0x0000040000400000) 
    12'hf58 : LOC <=          63'b000000000000000000001000000000000000000100000000000000000000000; // D (0x0000040000800000) 
    12'he8c : LOC <=          63'b000000000000000000001000000000000000001000000000000000000000000; // D (0x0000040001000000) 
    12'hd24 : LOC <=          63'b000000000000000000001000000000000000010000000000000000000000000; // D (0x0000040002000000) 
    12'ha74 : LOC <=          63'b000000000000000000001000000000000000100000000000000000000000000; // D (0x0000040004000000) 
    12'h4d4 : LOC <=          63'b000000000000000000001000000000000001000000000000000000000000000; // D (0x0000040008000000) 
    12'hcad : LOC <=          63'b000000000000000000001000000000000010000000000000000000000000000; // D (0x0000040010000000) 
    12'h966 : LOC <=          63'b000000000000000000001000000000000100000000000000000000000000000; // D (0x0000040020000000) 
    12'h2f0 : LOC <=          63'b000000000000000000001000000000001000000000000000000000000000000; // D (0x0000040040000000) 
    12'h0e5 : LOC <=          63'b000000000000000000001000000000010000000000000000000000000000000; // D (0x0000040080000000) 
    12'h4cf : LOC <=          63'b000000000000000000001000000000100000000000000000000000000000000; // D (0x0000040100000000) 
    12'hc9b : LOC <=          63'b000000000000000000001000000001000000000000000000000000000000000; // D (0x0000040200000000) 
    12'h90a : LOC <=          63'b000000000000000000001000000010000000000000000000000000000000000; // D (0x0000040400000000) 
    12'h228 : LOC <=          63'b000000000000000000001000000100000000000000000000000000000000000; // D (0x0000040800000000) 
    12'h155 : LOC <=          63'b000000000000000000001000001000000000000000000000000000000000000; // D (0x0000041000000000) 
    12'h7af : LOC <=          63'b000000000000000000001000010000000000000000000000000000000000000; // D (0x0000042000000000) 
    12'ha5b : LOC <=          63'b000000000000000000001000100000000000000000000000000000000000000; // D (0x0000044000000000) 
    12'h48a : LOC <=          63'b000000000000000000001001000000000000000000000000000000000000000; // D (0x0000048000000000) 
    12'hc11 : LOC <=          63'b000000000000000000001010000000000000000000000000000000000000000; // D (0x0000050000000000) 
    12'h81e : LOC <=          63'b000000000000000000001100000000000000000000000000000000000000000; // D (0x0000060000000000) 
    12'h303 : LOC <=          63'b000000000000000000001000000000000000000000000000000000000000000; // S (0x0000040000000000) 
//    12'h505 : LOC <=          63'b000000000000000000011000000000000000000000000000000000000000000; // D (0x00000c0000000000) 
//    12'hf0f : LOC <=          63'b000000000000000000101000000000000000000000000000000000000000000; // D (0x0000140000000000) 
//    12'he22 : LOC <=          63'b000000000000000001001000000000000000000000000000000000000000000; // D (0x0000240000000000) 
//    12'hc78 : LOC <=          63'b000000000000000010001000000000000000000000000000000000000000000; // D (0x0000440000000000) 
//    12'h8cc : LOC <=          63'b000000000000000100001000000000000000000000000000000000000000000; // D (0x0000840000000000) 
//    12'h1a4 : LOC <=          63'b000000000000001000001000000000000000000000000000000000000000000; // D (0x0001040000000000) 
//    12'h64d : LOC <=          63'b000000000000010000001000000000000000000000000000000000000000000; // D (0x0002040000000000) 
//    12'h99f : LOC <=          63'b000000000000100000001000000000000000000000000000000000000000000; // D (0x0004040000000000) 
//    12'h302 : LOC <=          63'b000000000001000000001000000000000000000000000000000000000000000; // D (0x0008040000000000) 
//    12'h301 : LOC <=          63'b000000000010000000001000000000000000000000000000000000000000000; // D (0x0010040000000000) 
//    12'h307 : LOC <=          63'b000000000100000000001000000000000000000000000000000000000000000; // D (0x0020040000000000) 
//    12'h30b : LOC <=          63'b000000001000000000001000000000000000000000000000000000000000000; // D (0x0040040000000000) 
//    12'h313 : LOC <=          63'b000000010000000000001000000000000000000000000000000000000000000; // D (0x0080040000000000) 
//    12'h323 : LOC <=          63'b000000100000000000001000000000000000000000000000000000000000000; // D (0x0100040000000000) 
//    12'h343 : LOC <=          63'b000001000000000000001000000000000000000000000000000000000000000; // D (0x0200040000000000) 
//    12'h383 : LOC <=          63'b000010000000000000001000000000000000000000000000000000000000000; // D (0x0400040000000000) 
//    12'h203 : LOC <=          63'b000100000000000000001000000000000000000000000000000000000000000; // D (0x0800040000000000) 
//    12'h103 : LOC <=          63'b001000000000000000001000000000000000000000000000000000000000000; // D (0x1000040000000000) 
//    12'h703 : LOC <=          63'b010000000000000000001000000000000000000000000000000000000000000; // D (0x2000040000000000) 
//    12'hb03 : LOC <=          63'b100000000000000000001000000000000000000000000000000000000000000; // D (0x4000040000000000) 
    12'h33f : LOC <=          63'b000000000000000000010000000000000000000000000000000000000000001; // D (0x0000080000000001) 
    12'hc74 : LOC <=          63'b000000000000000000010000000000000000000000000000000000000000010; // D (0x0000080000000002) 
    12'h7db : LOC <=          63'b000000000000000000010000000000000000000000000000000000000000100; // D (0x0000080000000004) 
    12'h5bc : LOC <=          63'b000000000000000000010000000000000000000000000000000000000001000; // D (0x0000080000000008) 
    12'h172 : LOC <=          63'b000000000000000000010000000000000000000000000000000000000010000; // D (0x0000080000000010) 
    12'h8ee : LOC <=          63'b000000000000000000010000000000000000000000000000000000000100000; // D (0x0000080000000020) 
    12'heef : LOC <=          63'b000000000000000000010000000000000000000000000000000000001000000; // D (0x0000080000000040) 
    12'h2ed : LOC <=          63'b000000000000000000010000000000000000000000000000000000010000000; // D (0x0000080000000080) 
    12'hfd0 : LOC <=          63'b000000000000000000010000000000000000000000000000000000100000000; // D (0x0000080000000100) 
    12'h093 : LOC <=          63'b000000000000000000010000000000000000000000000000000001000000000; // D (0x0000080000000200) 
    12'hb2c : LOC <=          63'b000000000000000000010000000000000000000000000000000010000000000; // D (0x0000080000000400) 
    12'h96b : LOC <=          63'b000000000000000000010000000000000000000000000000000100000000000; // D (0x0000080000000800) 
    12'hde5 : LOC <=          63'b000000000000000000010000000000000000000000000000001000000000000; // D (0x0000080000001000) 
    12'h4f9 : LOC <=          63'b000000000000000000010000000000000000000000000000010000000000000; // D (0x0000080000002000) 
    12'h3f8 : LOC <=          63'b000000000000000000010000000000000000000000000000100000000000000; // D (0x0000080000004000) 
    12'hdfa : LOC <=          63'b000000000000000000010000000000000000000000000001000000000000000; // D (0x0000080000008000) 
    12'h4c7 : LOC <=          63'b000000000000000000010000000000000000000000000010000000000000000; // D (0x0000080000010000) 
    12'h384 : LOC <=          63'b000000000000000000010000000000000000000000000100000000000000000; // D (0x0000080000020000) 
    12'hd02 : LOC <=          63'b000000000000000000010000000000000000000000001000000000000000000; // D (0x0000080000040000) 
    12'h537 : LOC <=          63'b000000000000000000010000000000000000000000010000000000000000000; // D (0x0000080000080000) 
    12'h064 : LOC <=          63'b000000000000000000010000000000000000000000100000000000000000000; // D (0x0000080000100000) 
    12'hac2 : LOC <=          63'b000000000000000000010000000000000000000001000000000000000000000; // D (0x0000080000200000) 
    12'hab7 : LOC <=          63'b000000000000000000010000000000000000000010000000000000000000000; // D (0x0000080000400000) 
    12'ha5d : LOC <=          63'b000000000000000000010000000000000000000100000000000000000000000; // D (0x0000080000800000) 
    12'hb89 : LOC <=          63'b000000000000000000010000000000000000001000000000000000000000000; // D (0x0000080001000000) 
    12'h821 : LOC <=          63'b000000000000000000010000000000000000010000000000000000000000000; // D (0x0000080002000000) 
    12'hf71 : LOC <=          63'b000000000000000000010000000000000000100000000000000000000000000; // D (0x0000080004000000) 
    12'h1d1 : LOC <=          63'b000000000000000000010000000000000001000000000000000000000000000; // D (0x0000080008000000) 
    12'h9a8 : LOC <=          63'b000000000000000000010000000000000010000000000000000000000000000; // D (0x0000080010000000) 
    12'hc63 : LOC <=          63'b000000000000000000010000000000000100000000000000000000000000000; // D (0x0000080020000000) 
    12'h7f5 : LOC <=          63'b000000000000000000010000000000001000000000000000000000000000000; // D (0x0000080040000000) 
    12'h5e0 : LOC <=          63'b000000000000000000010000000000010000000000000000000000000000000; // D (0x0000080080000000) 
    12'h1ca : LOC <=          63'b000000000000000000010000000000100000000000000000000000000000000; // D (0x0000080100000000) 
    12'h99e : LOC <=          63'b000000000000000000010000000001000000000000000000000000000000000; // D (0x0000080200000000) 
    12'hc0f : LOC <=          63'b000000000000000000010000000010000000000000000000000000000000000; // D (0x0000080400000000) 
    12'h72d : LOC <=          63'b000000000000000000010000000100000000000000000000000000000000000; // D (0x0000080800000000) 
    12'h450 : LOC <=          63'b000000000000000000010000001000000000000000000000000000000000000; // D (0x0000081000000000) 
    12'h2aa : LOC <=          63'b000000000000000000010000010000000000000000000000000000000000000; // D (0x0000082000000000) 
    12'hf5e : LOC <=          63'b000000000000000000010000100000000000000000000000000000000000000; // D (0x0000084000000000) 
    12'h18f : LOC <=          63'b000000000000000000010001000000000000000000000000000000000000000; // D (0x0000088000000000) 
    12'h914 : LOC <=          63'b000000000000000000010010000000000000000000000000000000000000000; // D (0x0000090000000000) 
    12'hd1b : LOC <=          63'b000000000000000000010100000000000000000000000000000000000000000; // D (0x00000a0000000000) 
    12'h505 : LOC <=          63'b000000000000000000011000000000000000000000000000000000000000000; // D (0x00000c0000000000) 
    12'h606 : LOC <=          63'b000000000000000000010000000000000000000000000000000000000000000; // S (0x0000080000000000) 
//    12'ha0a : LOC <=          63'b000000000000000000110000000000000000000000000000000000000000000; // D (0x0000180000000000) 
//    12'hb27 : LOC <=          63'b000000000000000001010000000000000000000000000000000000000000000; // D (0x0000280000000000) 
//    12'h97d : LOC <=          63'b000000000000000010010000000000000000000000000000000000000000000; // D (0x0000480000000000) 
//    12'hdc9 : LOC <=          63'b000000000000000100010000000000000000000000000000000000000000000; // D (0x0000880000000000) 
//    12'h4a1 : LOC <=          63'b000000000000001000010000000000000000000000000000000000000000000; // D (0x0001080000000000) 
//    12'h348 : LOC <=          63'b000000000000010000010000000000000000000000000000000000000000000; // D (0x0002080000000000) 
//    12'hc9a : LOC <=          63'b000000000000100000010000000000000000000000000000000000000000000; // D (0x0004080000000000) 
//    12'h607 : LOC <=          63'b000000000001000000010000000000000000000000000000000000000000000; // D (0x0008080000000000) 
//    12'h604 : LOC <=          63'b000000000010000000010000000000000000000000000000000000000000000; // D (0x0010080000000000) 
//    12'h602 : LOC <=          63'b000000000100000000010000000000000000000000000000000000000000000; // D (0x0020080000000000) 
//    12'h60e : LOC <=          63'b000000001000000000010000000000000000000000000000000000000000000; // D (0x0040080000000000) 
//    12'h616 : LOC <=          63'b000000010000000000010000000000000000000000000000000000000000000; // D (0x0080080000000000) 
//    12'h626 : LOC <=          63'b000000100000000000010000000000000000000000000000000000000000000; // D (0x0100080000000000) 
//    12'h646 : LOC <=          63'b000001000000000000010000000000000000000000000000000000000000000; // D (0x0200080000000000) 
//    12'h686 : LOC <=          63'b000010000000000000010000000000000000000000000000000000000000000; // D (0x0400080000000000) 
//    12'h706 : LOC <=          63'b000100000000000000010000000000000000000000000000000000000000000; // D (0x0800080000000000) 
//    12'h406 : LOC <=          63'b001000000000000000010000000000000000000000000000000000000000000; // D (0x1000080000000000) 
//    12'h206 : LOC <=          63'b010000000000000000010000000000000000000000000000000000000000000; // D (0x2000080000000000) 
//    12'he06 : LOC <=          63'b100000000000000000010000000000000000000000000000000000000000000; // D (0x4000080000000000) 
    12'h935 : LOC <=          63'b000000000000000000100000000000000000000000000000000000000000001; // D (0x0000100000000001) 
    12'h67e : LOC <=          63'b000000000000000000100000000000000000000000000000000000000000010; // D (0x0000100000000002) 
    12'hdd1 : LOC <=          63'b000000000000000000100000000000000000000000000000000000000000100; // D (0x0000100000000004) 
    12'hfb6 : LOC <=          63'b000000000000000000100000000000000000000000000000000000000001000; // D (0x0000100000000008) 
    12'hb78 : LOC <=          63'b000000000000000000100000000000000000000000000000000000000010000; // D (0x0000100000000010) 
    12'h2e4 : LOC <=          63'b000000000000000000100000000000000000000000000000000000000100000; // D (0x0000100000000020) 
    12'h4e5 : LOC <=          63'b000000000000000000100000000000000000000000000000000000001000000; // D (0x0000100000000040) 
    12'h8e7 : LOC <=          63'b000000000000000000100000000000000000000000000000000000010000000; // D (0x0000100000000080) 
    12'h5da : LOC <=          63'b000000000000000000100000000000000000000000000000000000100000000; // D (0x0000100000000100) 
    12'ha99 : LOC <=          63'b000000000000000000100000000000000000000000000000000001000000000; // D (0x0000100000000200) 
    12'h126 : LOC <=          63'b000000000000000000100000000000000000000000000000000010000000000; // D (0x0000100000000400) 
    12'h361 : LOC <=          63'b000000000000000000100000000000000000000000000000000100000000000; // D (0x0000100000000800) 
    12'h7ef : LOC <=          63'b000000000000000000100000000000000000000000000000001000000000000; // D (0x0000100000001000) 
    12'hef3 : LOC <=          63'b000000000000000000100000000000000000000000000000010000000000000; // D (0x0000100000002000) 
    12'h9f2 : LOC <=          63'b000000000000000000100000000000000000000000000000100000000000000; // D (0x0000100000004000) 
    12'h7f0 : LOC <=          63'b000000000000000000100000000000000000000000000001000000000000000; // D (0x0000100000008000) 
    12'hecd : LOC <=          63'b000000000000000000100000000000000000000000000010000000000000000; // D (0x0000100000010000) 
    12'h98e : LOC <=          63'b000000000000000000100000000000000000000000000100000000000000000; // D (0x0000100000020000) 
    12'h708 : LOC <=          63'b000000000000000000100000000000000000000000001000000000000000000; // D (0x0000100000040000) 
    12'hf3d : LOC <=          63'b000000000000000000100000000000000000000000010000000000000000000; // D (0x0000100000080000) 
    12'ha6e : LOC <=          63'b000000000000000000100000000000000000000000100000000000000000000; // D (0x0000100000100000) 
    12'h0c8 : LOC <=          63'b000000000000000000100000000000000000000001000000000000000000000; // D (0x0000100000200000) 
    12'h0bd : LOC <=          63'b000000000000000000100000000000000000000010000000000000000000000; // D (0x0000100000400000) 
    12'h057 : LOC <=          63'b000000000000000000100000000000000000000100000000000000000000000; // D (0x0000100000800000) 
    12'h183 : LOC <=          63'b000000000000000000100000000000000000001000000000000000000000000; // D (0x0000100001000000) 
    12'h22b : LOC <=          63'b000000000000000000100000000000000000010000000000000000000000000; // D (0x0000100002000000) 
    12'h57b : LOC <=          63'b000000000000000000100000000000000000100000000000000000000000000; // D (0x0000100004000000) 
    12'hbdb : LOC <=          63'b000000000000000000100000000000000001000000000000000000000000000; // D (0x0000100008000000) 
    12'h3a2 : LOC <=          63'b000000000000000000100000000000000010000000000000000000000000000; // D (0x0000100010000000) 
    12'h669 : LOC <=          63'b000000000000000000100000000000000100000000000000000000000000000; // D (0x0000100020000000) 
    12'hdff : LOC <=          63'b000000000000000000100000000000001000000000000000000000000000000; // D (0x0000100040000000) 
    12'hfea : LOC <=          63'b000000000000000000100000000000010000000000000000000000000000000; // D (0x0000100080000000) 
    12'hbc0 : LOC <=          63'b000000000000000000100000000000100000000000000000000000000000000; // D (0x0000100100000000) 
    12'h394 : LOC <=          63'b000000000000000000100000000001000000000000000000000000000000000; // D (0x0000100200000000) 
    12'h605 : LOC <=          63'b000000000000000000100000000010000000000000000000000000000000000; // D (0x0000100400000000) 
    12'hd27 : LOC <=          63'b000000000000000000100000000100000000000000000000000000000000000; // D (0x0000100800000000) 
    12'he5a : LOC <=          63'b000000000000000000100000001000000000000000000000000000000000000; // D (0x0000101000000000) 
    12'h8a0 : LOC <=          63'b000000000000000000100000010000000000000000000000000000000000000; // D (0x0000102000000000) 
    12'h554 : LOC <=          63'b000000000000000000100000100000000000000000000000000000000000000; // D (0x0000104000000000) 
    12'hb85 : LOC <=          63'b000000000000000000100001000000000000000000000000000000000000000; // D (0x0000108000000000) 
    12'h31e : LOC <=          63'b000000000000000000100010000000000000000000000000000000000000000; // D (0x0000110000000000) 
    12'h711 : LOC <=          63'b000000000000000000100100000000000000000000000000000000000000000; // D (0x0000120000000000) 
    12'hf0f : LOC <=          63'b000000000000000000101000000000000000000000000000000000000000000; // D (0x0000140000000000) 
    12'ha0a : LOC <=          63'b000000000000000000110000000000000000000000000000000000000000000; // D (0x0000180000000000) 
    12'hc0c : LOC <=          63'b000000000000000000100000000000000000000000000000000000000000000; // S (0x0000100000000000) 
//    12'h12d : LOC <=          63'b000000000000000001100000000000000000000000000000000000000000000; // D (0x0000300000000000) 
//    12'h377 : LOC <=          63'b000000000000000010100000000000000000000000000000000000000000000; // D (0x0000500000000000) 
//    12'h7c3 : LOC <=          63'b000000000000000100100000000000000000000000000000000000000000000; // D (0x0000900000000000) 
//    12'heab : LOC <=          63'b000000000000001000100000000000000000000000000000000000000000000; // D (0x0001100000000000) 
//    12'h942 : LOC <=          63'b000000000000010000100000000000000000000000000000000000000000000; // D (0x0002100000000000) 
//    12'h690 : LOC <=          63'b000000000000100000100000000000000000000000000000000000000000000; // D (0x0004100000000000) 
//    12'hc0d : LOC <=          63'b000000000001000000100000000000000000000000000000000000000000000; // D (0x0008100000000000) 
//    12'hc0e : LOC <=          63'b000000000010000000100000000000000000000000000000000000000000000; // D (0x0010100000000000) 
//    12'hc08 : LOC <=          63'b000000000100000000100000000000000000000000000000000000000000000; // D (0x0020100000000000) 
//    12'hc04 : LOC <=          63'b000000001000000000100000000000000000000000000000000000000000000; // D (0x0040100000000000) 
//    12'hc1c : LOC <=          63'b000000010000000000100000000000000000000000000000000000000000000; // D (0x0080100000000000) 
//    12'hc2c : LOC <=          63'b000000100000000000100000000000000000000000000000000000000000000; // D (0x0100100000000000) 
//    12'hc4c : LOC <=          63'b000001000000000000100000000000000000000000000000000000000000000; // D (0x0200100000000000) 
//    12'hc8c : LOC <=          63'b000010000000000000100000000000000000000000000000000000000000000; // D (0x0400100000000000) 
//    12'hd0c : LOC <=          63'b000100000000000000100000000000000000000000000000000000000000000; // D (0x0800100000000000) 
//    12'he0c : LOC <=          63'b001000000000000000100000000000000000000000000000000000000000000; // D (0x1000100000000000) 
//    12'h80c : LOC <=          63'b010000000000000000100000000000000000000000000000000000000000000; // D (0x2000100000000000) 
//    12'h40c : LOC <=          63'b100000000000000000100000000000000000000000000000000000000000000; // D (0x4000100000000000) 
    12'h818 : LOC <=          63'b000000000000000001000000000000000000000000000000000000000000001; // D (0x0000200000000001) 
    12'h753 : LOC <=          63'b000000000000000001000000000000000000000000000000000000000000010; // D (0x0000200000000002) 
    12'hcfc : LOC <=          63'b000000000000000001000000000000000000000000000000000000000000100; // D (0x0000200000000004) 
    12'he9b : LOC <=          63'b000000000000000001000000000000000000000000000000000000000001000; // D (0x0000200000000008) 
    12'ha55 : LOC <=          63'b000000000000000001000000000000000000000000000000000000000010000; // D (0x0000200000000010) 
    12'h3c9 : LOC <=          63'b000000000000000001000000000000000000000000000000000000000100000; // D (0x0000200000000020) 
    12'h5c8 : LOC <=          63'b000000000000000001000000000000000000000000000000000000001000000; // D (0x0000200000000040) 
    12'h9ca : LOC <=          63'b000000000000000001000000000000000000000000000000000000010000000; // D (0x0000200000000080) 
    12'h4f7 : LOC <=          63'b000000000000000001000000000000000000000000000000000000100000000; // D (0x0000200000000100) 
    12'hbb4 : LOC <=          63'b000000000000000001000000000000000000000000000000000001000000000; // D (0x0000200000000200) 
    12'h00b : LOC <=          63'b000000000000000001000000000000000000000000000000000010000000000; // D (0x0000200000000400) 
    12'h24c : LOC <=          63'b000000000000000001000000000000000000000000000000000100000000000; // D (0x0000200000000800) 
    12'h6c2 : LOC <=          63'b000000000000000001000000000000000000000000000000001000000000000; // D (0x0000200000001000) 
    12'hfde : LOC <=          63'b000000000000000001000000000000000000000000000000010000000000000; // D (0x0000200000002000) 
    12'h8df : LOC <=          63'b000000000000000001000000000000000000000000000000100000000000000; // D (0x0000200000004000) 
    12'h6dd : LOC <=          63'b000000000000000001000000000000000000000000000001000000000000000; // D (0x0000200000008000) 
    12'hfe0 : LOC <=          63'b000000000000000001000000000000000000000000000010000000000000000; // D (0x0000200000010000) 
    12'h8a3 : LOC <=          63'b000000000000000001000000000000000000000000000100000000000000000; // D (0x0000200000020000) 
    12'h625 : LOC <=          63'b000000000000000001000000000000000000000000001000000000000000000; // D (0x0000200000040000) 
    12'he10 : LOC <=          63'b000000000000000001000000000000000000000000010000000000000000000; // D (0x0000200000080000) 
    12'hb43 : LOC <=          63'b000000000000000001000000000000000000000000100000000000000000000; // D (0x0000200000100000) 
    12'h1e5 : LOC <=          63'b000000000000000001000000000000000000000001000000000000000000000; // D (0x0000200000200000) 
    12'h190 : LOC <=          63'b000000000000000001000000000000000000000010000000000000000000000; // D (0x0000200000400000) 
    12'h17a : LOC <=          63'b000000000000000001000000000000000000000100000000000000000000000; // D (0x0000200000800000) 
    12'h0ae : LOC <=          63'b000000000000000001000000000000000000001000000000000000000000000; // D (0x0000200001000000) 
    12'h306 : LOC <=          63'b000000000000000001000000000000000000010000000000000000000000000; // D (0x0000200002000000) 
    12'h456 : LOC <=          63'b000000000000000001000000000000000000100000000000000000000000000; // D (0x0000200004000000) 
    12'haf6 : LOC <=          63'b000000000000000001000000000000000001000000000000000000000000000; // D (0x0000200008000000) 
    12'h28f : LOC <=          63'b000000000000000001000000000000000010000000000000000000000000000; // D (0x0000200010000000) 
    12'h744 : LOC <=          63'b000000000000000001000000000000000100000000000000000000000000000; // D (0x0000200020000000) 
    12'hcd2 : LOC <=          63'b000000000000000001000000000000001000000000000000000000000000000; // D (0x0000200040000000) 
    12'hec7 : LOC <=          63'b000000000000000001000000000000010000000000000000000000000000000; // D (0x0000200080000000) 
    12'haed : LOC <=          63'b000000000000000001000000000000100000000000000000000000000000000; // D (0x0000200100000000) 
    12'h2b9 : LOC <=          63'b000000000000000001000000000001000000000000000000000000000000000; // D (0x0000200200000000) 
    12'h728 : LOC <=          63'b000000000000000001000000000010000000000000000000000000000000000; // D (0x0000200400000000) 
    12'hc0a : LOC <=          63'b000000000000000001000000000100000000000000000000000000000000000; // D (0x0000200800000000) 
    12'hf77 : LOC <=          63'b000000000000000001000000001000000000000000000000000000000000000; // D (0x0000201000000000) 
    12'h98d : LOC <=          63'b000000000000000001000000010000000000000000000000000000000000000; // D (0x0000202000000000) 
    12'h479 : LOC <=          63'b000000000000000001000000100000000000000000000000000000000000000; // D (0x0000204000000000) 
    12'haa8 : LOC <=          63'b000000000000000001000001000000000000000000000000000000000000000; // D (0x0000208000000000) 
    12'h233 : LOC <=          63'b000000000000000001000010000000000000000000000000000000000000000; // D (0x0000210000000000) 
    12'h63c : LOC <=          63'b000000000000000001000100000000000000000000000000000000000000000; // D (0x0000220000000000) 
    12'he22 : LOC <=          63'b000000000000000001001000000000000000000000000000000000000000000; // D (0x0000240000000000) 
    12'hb27 : LOC <=          63'b000000000000000001010000000000000000000000000000000000000000000; // D (0x0000280000000000) 
    12'h12d : LOC <=          63'b000000000000000001100000000000000000000000000000000000000000000; // D (0x0000300000000000) 
    12'hd21 : LOC <=          63'b000000000000000001000000000000000000000000000000000000000000000; // S (0x0000200000000000) 
//    12'h25a : LOC <=          63'b000000000000000011000000000000000000000000000000000000000000000; // D (0x0000600000000000) 
//    12'h6ee : LOC <=          63'b000000000000000101000000000000000000000000000000000000000000000; // D (0x0000a00000000000) 
//    12'hf86 : LOC <=          63'b000000000000001001000000000000000000000000000000000000000000000; // D (0x0001200000000000) 
//    12'h86f : LOC <=          63'b000000000000010001000000000000000000000000000000000000000000000; // D (0x0002200000000000) 
//    12'h7bd : LOC <=          63'b000000000000100001000000000000000000000000000000000000000000000; // D (0x0004200000000000) 
//    12'hd20 : LOC <=          63'b000000000001000001000000000000000000000000000000000000000000000; // D (0x0008200000000000) 
//    12'hd23 : LOC <=          63'b000000000010000001000000000000000000000000000000000000000000000; // D (0x0010200000000000) 
//    12'hd25 : LOC <=          63'b000000000100000001000000000000000000000000000000000000000000000; // D (0x0020200000000000) 
//    12'hd29 : LOC <=          63'b000000001000000001000000000000000000000000000000000000000000000; // D (0x0040200000000000) 
//    12'hd31 : LOC <=          63'b000000010000000001000000000000000000000000000000000000000000000; // D (0x0080200000000000) 
//    12'hd01 : LOC <=          63'b000000100000000001000000000000000000000000000000000000000000000; // D (0x0100200000000000) 
//    12'hd61 : LOC <=          63'b000001000000000001000000000000000000000000000000000000000000000; // D (0x0200200000000000) 
//    12'hda1 : LOC <=          63'b000010000000000001000000000000000000000000000000000000000000000; // D (0x0400200000000000) 
//    12'hc21 : LOC <=          63'b000100000000000001000000000000000000000000000000000000000000000; // D (0x0800200000000000) 
//    12'hf21 : LOC <=          63'b001000000000000001000000000000000000000000000000000000000000000; // D (0x1000200000000000) 
//    12'h921 : LOC <=          63'b010000000000000001000000000000000000000000000000000000000000000; // D (0x2000200000000000) 
//    12'h521 : LOC <=          63'b100000000000000001000000000000000000000000000000000000000000000; // D (0x4000200000000000) 
    12'ha42 : LOC <=          63'b000000000000000010000000000000000000000000000000000000000000001; // D (0x0000400000000001) 
    12'h509 : LOC <=          63'b000000000000000010000000000000000000000000000000000000000000010; // D (0x0000400000000002) 
    12'hea6 : LOC <=          63'b000000000000000010000000000000000000000000000000000000000000100; // D (0x0000400000000004) 
    12'hcc1 : LOC <=          63'b000000000000000010000000000000000000000000000000000000000001000; // D (0x0000400000000008) 
    12'h80f : LOC <=          63'b000000000000000010000000000000000000000000000000000000000010000; // D (0x0000400000000010) 
    12'h193 : LOC <=          63'b000000000000000010000000000000000000000000000000000000000100000; // D (0x0000400000000020) 
    12'h792 : LOC <=          63'b000000000000000010000000000000000000000000000000000000001000000; // D (0x0000400000000040) 
    12'hb90 : LOC <=          63'b000000000000000010000000000000000000000000000000000000010000000; // D (0x0000400000000080) 
    12'h6ad : LOC <=          63'b000000000000000010000000000000000000000000000000000000100000000; // D (0x0000400000000100) 
    12'h9ee : LOC <=          63'b000000000000000010000000000000000000000000000000000001000000000; // D (0x0000400000000200) 
    12'h251 : LOC <=          63'b000000000000000010000000000000000000000000000000000010000000000; // D (0x0000400000000400) 
    12'h016 : LOC <=          63'b000000000000000010000000000000000000000000000000000100000000000; // D (0x0000400000000800) 
    12'h498 : LOC <=          63'b000000000000000010000000000000000000000000000000001000000000000; // D (0x0000400000001000) 
    12'hd84 : LOC <=          63'b000000000000000010000000000000000000000000000000010000000000000; // D (0x0000400000002000) 
    12'ha85 : LOC <=          63'b000000000000000010000000000000000000000000000000100000000000000; // D (0x0000400000004000) 
    12'h487 : LOC <=          63'b000000000000000010000000000000000000000000000001000000000000000; // D (0x0000400000008000) 
    12'hdba : LOC <=          63'b000000000000000010000000000000000000000000000010000000000000000; // D (0x0000400000010000) 
    12'haf9 : LOC <=          63'b000000000000000010000000000000000000000000000100000000000000000; // D (0x0000400000020000) 
    12'h47f : LOC <=          63'b000000000000000010000000000000000000000000001000000000000000000; // D (0x0000400000040000) 
    12'hc4a : LOC <=          63'b000000000000000010000000000000000000000000010000000000000000000; // D (0x0000400000080000) 
    12'h919 : LOC <=          63'b000000000000000010000000000000000000000000100000000000000000000; // D (0x0000400000100000) 
    12'h3bf : LOC <=          63'b000000000000000010000000000000000000000001000000000000000000000; // D (0x0000400000200000) 
    12'h3ca : LOC <=          63'b000000000000000010000000000000000000000010000000000000000000000; // D (0x0000400000400000) 
    12'h320 : LOC <=          63'b000000000000000010000000000000000000000100000000000000000000000; // D (0x0000400000800000) 
    12'h2f4 : LOC <=          63'b000000000000000010000000000000000000001000000000000000000000000; // D (0x0000400001000000) 
    12'h15c : LOC <=          63'b000000000000000010000000000000000000010000000000000000000000000; // D (0x0000400002000000) 
    12'h60c : LOC <=          63'b000000000000000010000000000000000000100000000000000000000000000; // D (0x0000400004000000) 
    12'h8ac : LOC <=          63'b000000000000000010000000000000000001000000000000000000000000000; // D (0x0000400008000000) 
    12'h0d5 : LOC <=          63'b000000000000000010000000000000000010000000000000000000000000000; // D (0x0000400010000000) 
    12'h51e : LOC <=          63'b000000000000000010000000000000000100000000000000000000000000000; // D (0x0000400020000000) 
    12'he88 : LOC <=          63'b000000000000000010000000000000001000000000000000000000000000000; // D (0x0000400040000000) 
    12'hc9d : LOC <=          63'b000000000000000010000000000000010000000000000000000000000000000; // D (0x0000400080000000) 
    12'h8b7 : LOC <=          63'b000000000000000010000000000000100000000000000000000000000000000; // D (0x0000400100000000) 
    12'h0e3 : LOC <=          63'b000000000000000010000000000001000000000000000000000000000000000; // D (0x0000400200000000) 
    12'h572 : LOC <=          63'b000000000000000010000000000010000000000000000000000000000000000; // D (0x0000400400000000) 
    12'he50 : LOC <=          63'b000000000000000010000000000100000000000000000000000000000000000; // D (0x0000400800000000) 
    12'hd2d : LOC <=          63'b000000000000000010000000001000000000000000000000000000000000000; // D (0x0000401000000000) 
    12'hbd7 : LOC <=          63'b000000000000000010000000010000000000000000000000000000000000000; // D (0x0000402000000000) 
    12'h623 : LOC <=          63'b000000000000000010000000100000000000000000000000000000000000000; // D (0x0000404000000000) 
    12'h8f2 : LOC <=          63'b000000000000000010000001000000000000000000000000000000000000000; // D (0x0000408000000000) 
    12'h069 : LOC <=          63'b000000000000000010000010000000000000000000000000000000000000000; // D (0x0000410000000000) 
    12'h466 : LOC <=          63'b000000000000000010000100000000000000000000000000000000000000000; // D (0x0000420000000000) 
    12'hc78 : LOC <=          63'b000000000000000010001000000000000000000000000000000000000000000; // D (0x0000440000000000) 
    12'h97d : LOC <=          63'b000000000000000010010000000000000000000000000000000000000000000; // D (0x0000480000000000) 
    12'h377 : LOC <=          63'b000000000000000010100000000000000000000000000000000000000000000; // D (0x0000500000000000) 
    12'h25a : LOC <=          63'b000000000000000011000000000000000000000000000000000000000000000; // D (0x0000600000000000) 
    12'hf7b : LOC <=          63'b000000000000000010000000000000000000000000000000000000000000000; // S (0x0000400000000000) 
//    12'h4b4 : LOC <=          63'b000000000000000110000000000000000000000000000000000000000000000; // D (0x0000c00000000000) 
//    12'hddc : LOC <=          63'b000000000000001010000000000000000000000000000000000000000000000; // D (0x0001400000000000) 
//    12'ha35 : LOC <=          63'b000000000000010010000000000000000000000000000000000000000000000; // D (0x0002400000000000) 
//    12'h5e7 : LOC <=          63'b000000000000100010000000000000000000000000000000000000000000000; // D (0x0004400000000000) 
//    12'hf7a : LOC <=          63'b000000000001000010000000000000000000000000000000000000000000000; // D (0x0008400000000000) 
//    12'hf79 : LOC <=          63'b000000000010000010000000000000000000000000000000000000000000000; // D (0x0010400000000000) 
//    12'hf7f : LOC <=          63'b000000000100000010000000000000000000000000000000000000000000000; // D (0x0020400000000000) 
//    12'hf73 : LOC <=          63'b000000001000000010000000000000000000000000000000000000000000000; // D (0x0040400000000000) 
//    12'hf6b : LOC <=          63'b000000010000000010000000000000000000000000000000000000000000000; // D (0x0080400000000000) 
//    12'hf5b : LOC <=          63'b000000100000000010000000000000000000000000000000000000000000000; // D (0x0100400000000000) 
//    12'hf3b : LOC <=          63'b000001000000000010000000000000000000000000000000000000000000000; // D (0x0200400000000000) 
//    12'hffb : LOC <=          63'b000010000000000010000000000000000000000000000000000000000000000; // D (0x0400400000000000) 
//    12'he7b : LOC <=          63'b000100000000000010000000000000000000000000000000000000000000000; // D (0x0800400000000000) 
//    12'hd7b : LOC <=          63'b001000000000000010000000000000000000000000000000000000000000000; // D (0x1000400000000000) 
//    12'hb7b : LOC <=          63'b010000000000000010000000000000000000000000000000000000000000000; // D (0x2000400000000000) 
//    12'h77b : LOC <=          63'b100000000000000010000000000000000000000000000000000000000000000; // D (0x4000400000000000) 
    12'hef6 : LOC <=          63'b000000000000000100000000000000000000000000000000000000000000001; // D (0x0000800000000001) 
    12'h1bd : LOC <=          63'b000000000000000100000000000000000000000000000000000000000000010; // D (0x0000800000000002) 
    12'ha12 : LOC <=          63'b000000000000000100000000000000000000000000000000000000000000100; // D (0x0000800000000004) 
    12'h875 : LOC <=          63'b000000000000000100000000000000000000000000000000000000000001000; // D (0x0000800000000008) 
    12'hcbb : LOC <=          63'b000000000000000100000000000000000000000000000000000000000010000; // D (0x0000800000000010) 
    12'h527 : LOC <=          63'b000000000000000100000000000000000000000000000000000000000100000; // D (0x0000800000000020) 
    12'h326 : LOC <=          63'b000000000000000100000000000000000000000000000000000000001000000; // D (0x0000800000000040) 
    12'hf24 : LOC <=          63'b000000000000000100000000000000000000000000000000000000010000000; // D (0x0000800000000080) 
    12'h219 : LOC <=          63'b000000000000000100000000000000000000000000000000000000100000000; // D (0x0000800000000100) 
    12'hd5a : LOC <=          63'b000000000000000100000000000000000000000000000000000001000000000; // D (0x0000800000000200) 
    12'h6e5 : LOC <=          63'b000000000000000100000000000000000000000000000000000010000000000; // D (0x0000800000000400) 
    12'h4a2 : LOC <=          63'b000000000000000100000000000000000000000000000000000100000000000; // D (0x0000800000000800) 
    12'h02c : LOC <=          63'b000000000000000100000000000000000000000000000000001000000000000; // D (0x0000800000001000) 
    12'h930 : LOC <=          63'b000000000000000100000000000000000000000000000000010000000000000; // D (0x0000800000002000) 
    12'he31 : LOC <=          63'b000000000000000100000000000000000000000000000000100000000000000; // D (0x0000800000004000) 
    12'h033 : LOC <=          63'b000000000000000100000000000000000000000000000001000000000000000; // D (0x0000800000008000) 
    12'h90e : LOC <=          63'b000000000000000100000000000000000000000000000010000000000000000; // D (0x0000800000010000) 
    12'he4d : LOC <=          63'b000000000000000100000000000000000000000000000100000000000000000; // D (0x0000800000020000) 
    12'h0cb : LOC <=          63'b000000000000000100000000000000000000000000001000000000000000000; // D (0x0000800000040000) 
    12'h8fe : LOC <=          63'b000000000000000100000000000000000000000000010000000000000000000; // D (0x0000800000080000) 
    12'hdad : LOC <=          63'b000000000000000100000000000000000000000000100000000000000000000; // D (0x0000800000100000) 
    12'h70b : LOC <=          63'b000000000000000100000000000000000000000001000000000000000000000; // D (0x0000800000200000) 
    12'h77e : LOC <=          63'b000000000000000100000000000000000000000010000000000000000000000; // D (0x0000800000400000) 
    12'h794 : LOC <=          63'b000000000000000100000000000000000000000100000000000000000000000; // D (0x0000800000800000) 
    12'h640 : LOC <=          63'b000000000000000100000000000000000000001000000000000000000000000; // D (0x0000800001000000) 
    12'h5e8 : LOC <=          63'b000000000000000100000000000000000000010000000000000000000000000; // D (0x0000800002000000) 
    12'h2b8 : LOC <=          63'b000000000000000100000000000000000000100000000000000000000000000; // D (0x0000800004000000) 
    12'hc18 : LOC <=          63'b000000000000000100000000000000000001000000000000000000000000000; // D (0x0000800008000000) 
    12'h461 : LOC <=          63'b000000000000000100000000000000000010000000000000000000000000000; // D (0x0000800010000000) 
    12'h1aa : LOC <=          63'b000000000000000100000000000000000100000000000000000000000000000; // D (0x0000800020000000) 
    12'ha3c : LOC <=          63'b000000000000000100000000000000001000000000000000000000000000000; // D (0x0000800040000000) 
    12'h829 : LOC <=          63'b000000000000000100000000000000010000000000000000000000000000000; // D (0x0000800080000000) 
    12'hc03 : LOC <=          63'b000000000000000100000000000000100000000000000000000000000000000; // D (0x0000800100000000) 
    12'h457 : LOC <=          63'b000000000000000100000000000001000000000000000000000000000000000; // D (0x0000800200000000) 
    12'h1c6 : LOC <=          63'b000000000000000100000000000010000000000000000000000000000000000; // D (0x0000800400000000) 
    12'hae4 : LOC <=          63'b000000000000000100000000000100000000000000000000000000000000000; // D (0x0000800800000000) 
    12'h999 : LOC <=          63'b000000000000000100000000001000000000000000000000000000000000000; // D (0x0000801000000000) 
    12'hf63 : LOC <=          63'b000000000000000100000000010000000000000000000000000000000000000; // D (0x0000802000000000) 
    12'h297 : LOC <=          63'b000000000000000100000000100000000000000000000000000000000000000; // D (0x0000804000000000) 
    12'hc46 : LOC <=          63'b000000000000000100000001000000000000000000000000000000000000000; // D (0x0000808000000000) 
    12'h4dd : LOC <=          63'b000000000000000100000010000000000000000000000000000000000000000; // D (0x0000810000000000) 
    12'h0d2 : LOC <=          63'b000000000000000100000100000000000000000000000000000000000000000; // D (0x0000820000000000) 
    12'h8cc : LOC <=          63'b000000000000000100001000000000000000000000000000000000000000000; // D (0x0000840000000000) 
    12'hdc9 : LOC <=          63'b000000000000000100010000000000000000000000000000000000000000000; // D (0x0000880000000000) 
    12'h7c3 : LOC <=          63'b000000000000000100100000000000000000000000000000000000000000000; // D (0x0000900000000000) 
    12'h6ee : LOC <=          63'b000000000000000101000000000000000000000000000000000000000000000; // D (0x0000a00000000000) 
    12'h4b4 : LOC <=          63'b000000000000000110000000000000000000000000000000000000000000000; // D (0x0000c00000000000) 
    12'hbcf : LOC <=          63'b000000000000000100000000000000000000000000000000000000000000000; // S (0x0000800000000000) 
//    12'h968 : LOC <=          63'b000000000000001100000000000000000000000000000000000000000000000; // D (0x0001800000000000) 
//    12'he81 : LOC <=          63'b000000000000010100000000000000000000000000000000000000000000000; // D (0x0002800000000000) 
//    12'h153 : LOC <=          63'b000000000000100100000000000000000000000000000000000000000000000; // D (0x0004800000000000) 
//    12'hbce : LOC <=          63'b000000000001000100000000000000000000000000000000000000000000000; // D (0x0008800000000000) 
//    12'hbcd : LOC <=          63'b000000000010000100000000000000000000000000000000000000000000000; // D (0x0010800000000000) 
//    12'hbcb : LOC <=          63'b000000000100000100000000000000000000000000000000000000000000000; // D (0x0020800000000000) 
//    12'hbc7 : LOC <=          63'b000000001000000100000000000000000000000000000000000000000000000; // D (0x0040800000000000) 
//    12'hbdf : LOC <=          63'b000000010000000100000000000000000000000000000000000000000000000; // D (0x0080800000000000) 
//    12'hbef : LOC <=          63'b000000100000000100000000000000000000000000000000000000000000000; // D (0x0100800000000000) 
//    12'hb8f : LOC <=          63'b000001000000000100000000000000000000000000000000000000000000000; // D (0x0200800000000000) 
//    12'hb4f : LOC <=          63'b000010000000000100000000000000000000000000000000000000000000000; // D (0x0400800000000000) 
//    12'hacf : LOC <=          63'b000100000000000100000000000000000000000000000000000000000000000; // D (0x0800800000000000) 
//    12'h9cf : LOC <=          63'b001000000000000100000000000000000000000000000000000000000000000; // D (0x1000800000000000) 
//    12'hfcf : LOC <=          63'b010000000000000100000000000000000000000000000000000000000000000; // D (0x2000800000000000) 
//    12'h3cf : LOC <=          63'b100000000000000100000000000000000000000000000000000000000000000; // D (0x4000800000000000) 
    12'h79e : LOC <=          63'b000000000000001000000000000000000000000000000000000000000000001; // D (0x0001000000000001) 
    12'h8d5 : LOC <=          63'b000000000000001000000000000000000000000000000000000000000000010; // D (0x0001000000000002) 
    12'h37a : LOC <=          63'b000000000000001000000000000000000000000000000000000000000000100; // D (0x0001000000000004) 
    12'h11d : LOC <=          63'b000000000000001000000000000000000000000000000000000000000001000; // D (0x0001000000000008) 
    12'h5d3 : LOC <=          63'b000000000000001000000000000000000000000000000000000000000010000; // D (0x0001000000000010) 
    12'hc4f : LOC <=          63'b000000000000001000000000000000000000000000000000000000000100000; // D (0x0001000000000020) 
    12'ha4e : LOC <=          63'b000000000000001000000000000000000000000000000000000000001000000; // D (0x0001000000000040) 
    12'h64c : LOC <=          63'b000000000000001000000000000000000000000000000000000000010000000; // D (0x0001000000000080) 
    12'hb71 : LOC <=          63'b000000000000001000000000000000000000000000000000000000100000000; // D (0x0001000000000100) 
    12'h432 : LOC <=          63'b000000000000001000000000000000000000000000000000000001000000000; // D (0x0001000000000200) 
    12'hf8d : LOC <=          63'b000000000000001000000000000000000000000000000000000010000000000; // D (0x0001000000000400) 
    12'hdca : LOC <=          63'b000000000000001000000000000000000000000000000000000100000000000; // D (0x0001000000000800) 
    12'h944 : LOC <=          63'b000000000000001000000000000000000000000000000000001000000000000; // D (0x0001000000001000) 
    12'h058 : LOC <=          63'b000000000000001000000000000000000000000000000000010000000000000; // D (0x0001000000002000) 
    12'h759 : LOC <=          63'b000000000000001000000000000000000000000000000000100000000000000; // D (0x0001000000004000) 
    12'h95b : LOC <=          63'b000000000000001000000000000000000000000000000001000000000000000; // D (0x0001000000008000) 
    12'h066 : LOC <=          63'b000000000000001000000000000000000000000000000010000000000000000; // D (0x0001000000010000) 
    12'h725 : LOC <=          63'b000000000000001000000000000000000000000000000100000000000000000; // D (0x0001000000020000) 
    12'h9a3 : LOC <=          63'b000000000000001000000000000000000000000000001000000000000000000; // D (0x0001000000040000) 
    12'h196 : LOC <=          63'b000000000000001000000000000000000000000000010000000000000000000; // D (0x0001000000080000) 
    12'h4c5 : LOC <=          63'b000000000000001000000000000000000000000000100000000000000000000; // D (0x0001000000100000) 
    12'he63 : LOC <=          63'b000000000000001000000000000000000000000001000000000000000000000; // D (0x0001000000200000) 
    12'he16 : LOC <=          63'b000000000000001000000000000000000000000010000000000000000000000; // D (0x0001000000400000) 
    12'hefc : LOC <=          63'b000000000000001000000000000000000000000100000000000000000000000; // D (0x0001000000800000) 
    12'hf28 : LOC <=          63'b000000000000001000000000000000000000001000000000000000000000000; // D (0x0001000001000000) 
    12'hc80 : LOC <=          63'b000000000000001000000000000000000000010000000000000000000000000; // D (0x0001000002000000) 
    12'hbd0 : LOC <=          63'b000000000000001000000000000000000000100000000000000000000000000; // D (0x0001000004000000) 
    12'h570 : LOC <=          63'b000000000000001000000000000000000001000000000000000000000000000; // D (0x0001000008000000) 
    12'hd09 : LOC <=          63'b000000000000001000000000000000000010000000000000000000000000000; // D (0x0001000010000000) 
    12'h8c2 : LOC <=          63'b000000000000001000000000000000000100000000000000000000000000000; // D (0x0001000020000000) 
    12'h354 : LOC <=          63'b000000000000001000000000000000001000000000000000000000000000000; // D (0x0001000040000000) 
    12'h141 : LOC <=          63'b000000000000001000000000000000010000000000000000000000000000000; // D (0x0001000080000000) 
    12'h56b : LOC <=          63'b000000000000001000000000000000100000000000000000000000000000000; // D (0x0001000100000000) 
    12'hd3f : LOC <=          63'b000000000000001000000000000001000000000000000000000000000000000; // D (0x0001000200000000) 
    12'h8ae : LOC <=          63'b000000000000001000000000000010000000000000000000000000000000000; // D (0x0001000400000000) 
    12'h38c : LOC <=          63'b000000000000001000000000000100000000000000000000000000000000000; // D (0x0001000800000000) 
    12'h0f1 : LOC <=          63'b000000000000001000000000001000000000000000000000000000000000000; // D (0x0001001000000000) 
    12'h60b : LOC <=          63'b000000000000001000000000010000000000000000000000000000000000000; // D (0x0001002000000000) 
    12'hbff : LOC <=          63'b000000000000001000000000100000000000000000000000000000000000000; // D (0x0001004000000000) 
    12'h52e : LOC <=          63'b000000000000001000000001000000000000000000000000000000000000000; // D (0x0001008000000000) 
    12'hdb5 : LOC <=          63'b000000000000001000000010000000000000000000000000000000000000000; // D (0x0001010000000000) 
    12'h9ba : LOC <=          63'b000000000000001000000100000000000000000000000000000000000000000; // D (0x0001020000000000) 
    12'h1a4 : LOC <=          63'b000000000000001000001000000000000000000000000000000000000000000; // D (0x0001040000000000) 
    12'h4a1 : LOC <=          63'b000000000000001000010000000000000000000000000000000000000000000; // D (0x0001080000000000) 
    12'heab : LOC <=          63'b000000000000001000100000000000000000000000000000000000000000000; // D (0x0001100000000000) 
    12'hf86 : LOC <=          63'b000000000000001001000000000000000000000000000000000000000000000; // D (0x0001200000000000) 
    12'hddc : LOC <=          63'b000000000000001010000000000000000000000000000000000000000000000; // D (0x0001400000000000) 
    12'h968 : LOC <=          63'b000000000000001100000000000000000000000000000000000000000000000; // D (0x0001800000000000) 
    12'h2a7 : LOC <=          63'b000000000000001000000000000000000000000000000000000000000000000; // S (0x0001000000000000) 
//    12'h7e9 : LOC <=          63'b000000000000011000000000000000000000000000000000000000000000000; // D (0x0003000000000000) 
//    12'h83b : LOC <=          63'b000000000000101000000000000000000000000000000000000000000000000; // D (0x0005000000000000) 
//    12'h2a6 : LOC <=          63'b000000000001001000000000000000000000000000000000000000000000000; // D (0x0009000000000000) 
//    12'h2a5 : LOC <=          63'b000000000010001000000000000000000000000000000000000000000000000; // D (0x0011000000000000) 
//    12'h2a3 : LOC <=          63'b000000000100001000000000000000000000000000000000000000000000000; // D (0x0021000000000000) 
//    12'h2af : LOC <=          63'b000000001000001000000000000000000000000000000000000000000000000; // D (0x0041000000000000) 
//    12'h2b7 : LOC <=          63'b000000010000001000000000000000000000000000000000000000000000000; // D (0x0081000000000000) 
//    12'h287 : LOC <=          63'b000000100000001000000000000000000000000000000000000000000000000; // D (0x0101000000000000) 
//    12'h2e7 : LOC <=          63'b000001000000001000000000000000000000000000000000000000000000000; // D (0x0201000000000000) 
//    12'h227 : LOC <=          63'b000010000000001000000000000000000000000000000000000000000000000; // D (0x0401000000000000) 
//    12'h3a7 : LOC <=          63'b000100000000001000000000000000000000000000000000000000000000000; // D (0x0801000000000000) 
//    12'h0a7 : LOC <=          63'b001000000000001000000000000000000000000000000000000000000000000; // D (0x1001000000000000) 
//    12'h6a7 : LOC <=          63'b010000000000001000000000000000000000000000000000000000000000000; // D (0x2001000000000000) 
//    12'haa7 : LOC <=          63'b100000000000001000000000000000000000000000000000000000000000000; // D (0x4001000000000000) 
    12'h077 : LOC <=          63'b000000000000010000000000000000000000000000000000000000000000001; // D (0x0002000000000001) 
    12'hf3c : LOC <=          63'b000000000000010000000000000000000000000000000000000000000000010; // D (0x0002000000000002) 
    12'h493 : LOC <=          63'b000000000000010000000000000000000000000000000000000000000000100; // D (0x0002000000000004) 
    12'h6f4 : LOC <=          63'b000000000000010000000000000000000000000000000000000000000001000; // D (0x0002000000000008) 
    12'h23a : LOC <=          63'b000000000000010000000000000000000000000000000000000000000010000; // D (0x0002000000000010) 
    12'hba6 : LOC <=          63'b000000000000010000000000000000000000000000000000000000000100000; // D (0x0002000000000020) 
    12'hda7 : LOC <=          63'b000000000000010000000000000000000000000000000000000000001000000; // D (0x0002000000000040) 
    12'h1a5 : LOC <=          63'b000000000000010000000000000000000000000000000000000000010000000; // D (0x0002000000000080) 
    12'hc98 : LOC <=          63'b000000000000010000000000000000000000000000000000000000100000000; // D (0x0002000000000100) 
    12'h3db : LOC <=          63'b000000000000010000000000000000000000000000000000000001000000000; // D (0x0002000000000200) 
    12'h864 : LOC <=          63'b000000000000010000000000000000000000000000000000000010000000000; // D (0x0002000000000400) 
    12'ha23 : LOC <=          63'b000000000000010000000000000000000000000000000000000100000000000; // D (0x0002000000000800) 
    12'head : LOC <=          63'b000000000000010000000000000000000000000000000000001000000000000; // D (0x0002000000001000) 
    12'h7b1 : LOC <=          63'b000000000000010000000000000000000000000000000000010000000000000; // D (0x0002000000002000) 
    12'h0b0 : LOC <=          63'b000000000000010000000000000000000000000000000000100000000000000; // D (0x0002000000004000) 
    12'heb2 : LOC <=          63'b000000000000010000000000000000000000000000000001000000000000000; // D (0x0002000000008000) 
    12'h78f : LOC <=          63'b000000000000010000000000000000000000000000000010000000000000000; // D (0x0002000000010000) 
    12'h0cc : LOC <=          63'b000000000000010000000000000000000000000000000100000000000000000; // D (0x0002000000020000) 
    12'he4a : LOC <=          63'b000000000000010000000000000000000000000000001000000000000000000; // D (0x0002000000040000) 
    12'h67f : LOC <=          63'b000000000000010000000000000000000000000000010000000000000000000; // D (0x0002000000080000) 
    12'h32c : LOC <=          63'b000000000000010000000000000000000000000000100000000000000000000; // D (0x0002000000100000) 
    12'h98a : LOC <=          63'b000000000000010000000000000000000000000001000000000000000000000; // D (0x0002000000200000) 
    12'h9ff : LOC <=          63'b000000000000010000000000000000000000000010000000000000000000000; // D (0x0002000000400000) 
    12'h915 : LOC <=          63'b000000000000010000000000000000000000000100000000000000000000000; // D (0x0002000000800000) 
    12'h8c1 : LOC <=          63'b000000000000010000000000000000000000001000000000000000000000000; // D (0x0002000001000000) 
    12'hb69 : LOC <=          63'b000000000000010000000000000000000000010000000000000000000000000; // D (0x0002000002000000) 
    12'hc39 : LOC <=          63'b000000000000010000000000000000000000100000000000000000000000000; // D (0x0002000004000000) 
    12'h299 : LOC <=          63'b000000000000010000000000000000000001000000000000000000000000000; // D (0x0002000008000000) 
    12'hae0 : LOC <=          63'b000000000000010000000000000000000010000000000000000000000000000; // D (0x0002000010000000) 
    12'hf2b : LOC <=          63'b000000000000010000000000000000000100000000000000000000000000000; // D (0x0002000020000000) 
    12'h4bd : LOC <=          63'b000000000000010000000000000000001000000000000000000000000000000; // D (0x0002000040000000) 
    12'h6a8 : LOC <=          63'b000000000000010000000000000000010000000000000000000000000000000; // D (0x0002000080000000) 
    12'h282 : LOC <=          63'b000000000000010000000000000000100000000000000000000000000000000; // D (0x0002000100000000) 
    12'had6 : LOC <=          63'b000000000000010000000000000001000000000000000000000000000000000; // D (0x0002000200000000) 
    12'hf47 : LOC <=          63'b000000000000010000000000000010000000000000000000000000000000000; // D (0x0002000400000000) 
    12'h465 : LOC <=          63'b000000000000010000000000000100000000000000000000000000000000000; // D (0x0002000800000000) 
    12'h718 : LOC <=          63'b000000000000010000000000001000000000000000000000000000000000000; // D (0x0002001000000000) 
    12'h1e2 : LOC <=          63'b000000000000010000000000010000000000000000000000000000000000000; // D (0x0002002000000000) 
    12'hc16 : LOC <=          63'b000000000000010000000000100000000000000000000000000000000000000; // D (0x0002004000000000) 
    12'h2c7 : LOC <=          63'b000000000000010000000001000000000000000000000000000000000000000; // D (0x0002008000000000) 
    12'ha5c : LOC <=          63'b000000000000010000000010000000000000000000000000000000000000000; // D (0x0002010000000000) 
    12'he53 : LOC <=          63'b000000000000010000000100000000000000000000000000000000000000000; // D (0x0002020000000000) 
    12'h64d : LOC <=          63'b000000000000010000001000000000000000000000000000000000000000000; // D (0x0002040000000000) 
    12'h348 : LOC <=          63'b000000000000010000010000000000000000000000000000000000000000000; // D (0x0002080000000000) 
    12'h942 : LOC <=          63'b000000000000010000100000000000000000000000000000000000000000000; // D (0x0002100000000000) 
    12'h86f : LOC <=          63'b000000000000010001000000000000000000000000000000000000000000000; // D (0x0002200000000000) 
    12'ha35 : LOC <=          63'b000000000000010010000000000000000000000000000000000000000000000; // D (0x0002400000000000) 
    12'he81 : LOC <=          63'b000000000000010100000000000000000000000000000000000000000000000; // D (0x0002800000000000) 
    12'h7e9 : LOC <=          63'b000000000000011000000000000000000000000000000000000000000000000; // D (0x0003000000000000) 
    12'h54e : LOC <=          63'b000000000000010000000000000000000000000000000000000000000000000; // S (0x0002000000000000) 
//    12'hfd2 : LOC <=          63'b000000000000110000000000000000000000000000000000000000000000000; // D (0x0006000000000000) 
//    12'h54f : LOC <=          63'b000000000001010000000000000000000000000000000000000000000000000; // D (0x000a000000000000) 
//    12'h54c : LOC <=          63'b000000000010010000000000000000000000000000000000000000000000000; // D (0x0012000000000000) 
//    12'h54a : LOC <=          63'b000000000100010000000000000000000000000000000000000000000000000; // D (0x0022000000000000) 
//    12'h546 : LOC <=          63'b000000001000010000000000000000000000000000000000000000000000000; // D (0x0042000000000000) 
//    12'h55e : LOC <=          63'b000000010000010000000000000000000000000000000000000000000000000; // D (0x0082000000000000) 
//    12'h56e : LOC <=          63'b000000100000010000000000000000000000000000000000000000000000000; // D (0x0102000000000000) 
//    12'h50e : LOC <=          63'b000001000000010000000000000000000000000000000000000000000000000; // D (0x0202000000000000) 
//    12'h5ce : LOC <=          63'b000010000000010000000000000000000000000000000000000000000000000; // D (0x0402000000000000) 
//    12'h44e : LOC <=          63'b000100000000010000000000000000000000000000000000000000000000000; // D (0x0802000000000000) 
//    12'h74e : LOC <=          63'b001000000000010000000000000000000000000000000000000000000000000; // D (0x1002000000000000) 
//    12'h14e : LOC <=          63'b010000000000010000000000000000000000000000000000000000000000000; // D (0x2002000000000000) 
//    12'hd4e : LOC <=          63'b100000000000010000000000000000000000000000000000000000000000000; // D (0x4002000000000000) 
    12'hfa5 : LOC <=          63'b000000000000100000000000000000000000000000000000000000000000001; // D (0x0004000000000001) 
    12'h0ee : LOC <=          63'b000000000000100000000000000000000000000000000000000000000000010; // D (0x0004000000000002) 
    12'hb41 : LOC <=          63'b000000000000100000000000000000000000000000000000000000000000100; // D (0x0004000000000004) 
    12'h926 : LOC <=          63'b000000000000100000000000000000000000000000000000000000000001000; // D (0x0004000000000008) 
    12'hde8 : LOC <=          63'b000000000000100000000000000000000000000000000000000000000010000; // D (0x0004000000000010) 
    12'h474 : LOC <=          63'b000000000000100000000000000000000000000000000000000000000100000; // D (0x0004000000000020) 
    12'h275 : LOC <=          63'b000000000000100000000000000000000000000000000000000000001000000; // D (0x0004000000000040) 
    12'he77 : LOC <=          63'b000000000000100000000000000000000000000000000000000000010000000; // D (0x0004000000000080) 
    12'h34a : LOC <=          63'b000000000000100000000000000000000000000000000000000000100000000; // D (0x0004000000000100) 
    12'hc09 : LOC <=          63'b000000000000100000000000000000000000000000000000000001000000000; // D (0x0004000000000200) 
    12'h7b6 : LOC <=          63'b000000000000100000000000000000000000000000000000000010000000000; // D (0x0004000000000400) 
    12'h5f1 : LOC <=          63'b000000000000100000000000000000000000000000000000000100000000000; // D (0x0004000000000800) 
    12'h17f : LOC <=          63'b000000000000100000000000000000000000000000000000001000000000000; // D (0x0004000000001000) 
    12'h863 : LOC <=          63'b000000000000100000000000000000000000000000000000010000000000000; // D (0x0004000000002000) 
    12'hf62 : LOC <=          63'b000000000000100000000000000000000000000000000000100000000000000; // D (0x0004000000004000) 
    12'h160 : LOC <=          63'b000000000000100000000000000000000000000000000001000000000000000; // D (0x0004000000008000) 
    12'h85d : LOC <=          63'b000000000000100000000000000000000000000000000010000000000000000; // D (0x0004000000010000) 
    12'hf1e : LOC <=          63'b000000000000100000000000000000000000000000000100000000000000000; // D (0x0004000000020000) 
    12'h198 : LOC <=          63'b000000000000100000000000000000000000000000001000000000000000000; // D (0x0004000000040000) 
    12'h9ad : LOC <=          63'b000000000000100000000000000000000000000000010000000000000000000; // D (0x0004000000080000) 
    12'hcfe : LOC <=          63'b000000000000100000000000000000000000000000100000000000000000000; // D (0x0004000000100000) 
    12'h658 : LOC <=          63'b000000000000100000000000000000000000000001000000000000000000000; // D (0x0004000000200000) 
    12'h62d : LOC <=          63'b000000000000100000000000000000000000000010000000000000000000000; // D (0x0004000000400000) 
    12'h6c7 : LOC <=          63'b000000000000100000000000000000000000000100000000000000000000000; // D (0x0004000000800000) 
    12'h713 : LOC <=          63'b000000000000100000000000000000000000001000000000000000000000000; // D (0x0004000001000000) 
    12'h4bb : LOC <=          63'b000000000000100000000000000000000000010000000000000000000000000; // D (0x0004000002000000) 
    12'h3eb : LOC <=          63'b000000000000100000000000000000000000100000000000000000000000000; // D (0x0004000004000000) 
    12'hd4b : LOC <=          63'b000000000000100000000000000000000001000000000000000000000000000; // D (0x0004000008000000) 
    12'h532 : LOC <=          63'b000000000000100000000000000000000010000000000000000000000000000; // D (0x0004000010000000) 
    12'h0f9 : LOC <=          63'b000000000000100000000000000000000100000000000000000000000000000; // D (0x0004000020000000) 
    12'hb6f : LOC <=          63'b000000000000100000000000000000001000000000000000000000000000000; // D (0x0004000040000000) 
    12'h97a : LOC <=          63'b000000000000100000000000000000010000000000000000000000000000000; // D (0x0004000080000000) 
    12'hd50 : LOC <=          63'b000000000000100000000000000000100000000000000000000000000000000; // D (0x0004000100000000) 
    12'h504 : LOC <=          63'b000000000000100000000000000001000000000000000000000000000000000; // D (0x0004000200000000) 
    12'h095 : LOC <=          63'b000000000000100000000000000010000000000000000000000000000000000; // D (0x0004000400000000) 
    12'hbb7 : LOC <=          63'b000000000000100000000000000100000000000000000000000000000000000; // D (0x0004000800000000) 
    12'h8ca : LOC <=          63'b000000000000100000000000001000000000000000000000000000000000000; // D (0x0004001000000000) 
    12'he30 : LOC <=          63'b000000000000100000000000010000000000000000000000000000000000000; // D (0x0004002000000000) 
    12'h3c4 : LOC <=          63'b000000000000100000000000100000000000000000000000000000000000000; // D (0x0004004000000000) 
    12'hd15 : LOC <=          63'b000000000000100000000001000000000000000000000000000000000000000; // D (0x0004008000000000) 
    12'h58e : LOC <=          63'b000000000000100000000010000000000000000000000000000000000000000; // D (0x0004010000000000) 
    12'h181 : LOC <=          63'b000000000000100000000100000000000000000000000000000000000000000; // D (0x0004020000000000) 
    12'h99f : LOC <=          63'b000000000000100000001000000000000000000000000000000000000000000; // D (0x0004040000000000) 
    12'hc9a : LOC <=          63'b000000000000100000010000000000000000000000000000000000000000000; // D (0x0004080000000000) 
    12'h690 : LOC <=          63'b000000000000100000100000000000000000000000000000000000000000000; // D (0x0004100000000000) 
    12'h7bd : LOC <=          63'b000000000000100001000000000000000000000000000000000000000000000; // D (0x0004200000000000) 
    12'h5e7 : LOC <=          63'b000000000000100010000000000000000000000000000000000000000000000; // D (0x0004400000000000) 
    12'h153 : LOC <=          63'b000000000000100100000000000000000000000000000000000000000000000; // D (0x0004800000000000) 
    12'h83b : LOC <=          63'b000000000000101000000000000000000000000000000000000000000000000; // D (0x0005000000000000) 
    12'hfd2 : LOC <=          63'b000000000000110000000000000000000000000000000000000000000000000; // D (0x0006000000000000) 
    12'ha9c : LOC <=          63'b000000000000100000000000000000000000000000000000000000000000000; // S (0x0004000000000000) 
//    12'ha9d : LOC <=          63'b000000000001100000000000000000000000000000000000000000000000000; // D (0x000c000000000000) 
//    12'ha9e : LOC <=          63'b000000000010100000000000000000000000000000000000000000000000000; // D (0x0014000000000000) 
//    12'ha98 : LOC <=          63'b000000000100100000000000000000000000000000000000000000000000000; // D (0x0024000000000000) 
//    12'ha94 : LOC <=          63'b000000001000100000000000000000000000000000000000000000000000000; // D (0x0044000000000000) 
//    12'ha8c : LOC <=          63'b000000010000100000000000000000000000000000000000000000000000000; // D (0x0084000000000000) 
//    12'habc : LOC <=          63'b000000100000100000000000000000000000000000000000000000000000000; // D (0x0104000000000000) 
//    12'hadc : LOC <=          63'b000001000000100000000000000000000000000000000000000000000000000; // D (0x0204000000000000) 
//    12'ha1c : LOC <=          63'b000010000000100000000000000000000000000000000000000000000000000; // D (0x0404000000000000) 
//    12'hb9c : LOC <=          63'b000100000000100000000000000000000000000000000000000000000000000; // D (0x0804000000000000) 
//    12'h89c : LOC <=          63'b001000000000100000000000000000000000000000000000000000000000000; // D (0x1004000000000000) 
//    12'he9c : LOC <=          63'b010000000000100000000000000000000000000000000000000000000000000; // D (0x2004000000000000) 
//    12'h29c : LOC <=          63'b100000000000100000000000000000000000000000000000000000000000000; // D (0x4004000000000000) 
    12'h538 : LOC <=          63'b000000000001000000000000000000000000000000000000000000000000001; // D (0x0008000000000001) 
    12'ha73 : LOC <=          63'b000000000001000000000000000000000000000000000000000000000000010; // D (0x0008000000000002) 
    12'h1dc : LOC <=          63'b000000000001000000000000000000000000000000000000000000000000100; // D (0x0008000000000004) 
    12'h3bb : LOC <=          63'b000000000001000000000000000000000000000000000000000000000001000; // D (0x0008000000000008) 
    12'h775 : LOC <=          63'b000000000001000000000000000000000000000000000000000000000010000; // D (0x0008000000000010) 
    12'hee9 : LOC <=          63'b000000000001000000000000000000000000000000000000000000000100000; // D (0x0008000000000020) 
    12'h8e8 : LOC <=          63'b000000000001000000000000000000000000000000000000000000001000000; // D (0x0008000000000040) 
    12'h4ea : LOC <=          63'b000000000001000000000000000000000000000000000000000000010000000; // D (0x0008000000000080) 
    12'h9d7 : LOC <=          63'b000000000001000000000000000000000000000000000000000000100000000; // D (0x0008000000000100) 
    12'h694 : LOC <=          63'b000000000001000000000000000000000000000000000000000001000000000; // D (0x0008000000000200) 
    12'hd2b : LOC <=          63'b000000000001000000000000000000000000000000000000000010000000000; // D (0x0008000000000400) 
    12'hf6c : LOC <=          63'b000000000001000000000000000000000000000000000000000100000000000; // D (0x0008000000000800) 
    12'hbe2 : LOC <=          63'b000000000001000000000000000000000000000000000000001000000000000; // D (0x0008000000001000) 
    12'h2fe : LOC <=          63'b000000000001000000000000000000000000000000000000010000000000000; // D (0x0008000000002000) 
    12'h5ff : LOC <=          63'b000000000001000000000000000000000000000000000000100000000000000; // D (0x0008000000004000) 
    12'hbfd : LOC <=          63'b000000000001000000000000000000000000000000000001000000000000000; // D (0x0008000000008000) 
    12'h2c0 : LOC <=          63'b000000000001000000000000000000000000000000000010000000000000000; // D (0x0008000000010000) 
    12'h583 : LOC <=          63'b000000000001000000000000000000000000000000000100000000000000000; // D (0x0008000000020000) 
    12'hb05 : LOC <=          63'b000000000001000000000000000000000000000000001000000000000000000; // D (0x0008000000040000) 
    12'h330 : LOC <=          63'b000000000001000000000000000000000000000000010000000000000000000; // D (0x0008000000080000) 
    12'h663 : LOC <=          63'b000000000001000000000000000000000000000000100000000000000000000; // D (0x0008000000100000) 
    12'hcc5 : LOC <=          63'b000000000001000000000000000000000000000001000000000000000000000; // D (0x0008000000200000) 
    12'hcb0 : LOC <=          63'b000000000001000000000000000000000000000010000000000000000000000; // D (0x0008000000400000) 
    12'hc5a : LOC <=          63'b000000000001000000000000000000000000000100000000000000000000000; // D (0x0008000000800000) 
    12'hd8e : LOC <=          63'b000000000001000000000000000000000000001000000000000000000000000; // D (0x0008000001000000) 
    12'he26 : LOC <=          63'b000000000001000000000000000000000000010000000000000000000000000; // D (0x0008000002000000) 
    12'h976 : LOC <=          63'b000000000001000000000000000000000000100000000000000000000000000; // D (0x0008000004000000) 
    12'h7d6 : LOC <=          63'b000000000001000000000000000000000001000000000000000000000000000; // D (0x0008000008000000) 
    12'hfaf : LOC <=          63'b000000000001000000000000000000000010000000000000000000000000000; // D (0x0008000010000000) 
    12'ha64 : LOC <=          63'b000000000001000000000000000000000100000000000000000000000000000; // D (0x0008000020000000) 
    12'h1f2 : LOC <=          63'b000000000001000000000000000000001000000000000000000000000000000; // D (0x0008000040000000) 
    12'h3e7 : LOC <=          63'b000000000001000000000000000000010000000000000000000000000000000; // D (0x0008000080000000) 
    12'h7cd : LOC <=          63'b000000000001000000000000000000100000000000000000000000000000000; // D (0x0008000100000000) 
    12'hf99 : LOC <=          63'b000000000001000000000000000001000000000000000000000000000000000; // D (0x0008000200000000) 
    12'ha08 : LOC <=          63'b000000000001000000000000000010000000000000000000000000000000000; // D (0x0008000400000000) 
    12'h12a : LOC <=          63'b000000000001000000000000000100000000000000000000000000000000000; // D (0x0008000800000000) 
    12'h257 : LOC <=          63'b000000000001000000000000001000000000000000000000000000000000000; // D (0x0008001000000000) 
    12'h4ad : LOC <=          63'b000000000001000000000000010000000000000000000000000000000000000; // D (0x0008002000000000) 
    12'h959 : LOC <=          63'b000000000001000000000000100000000000000000000000000000000000000; // D (0x0008004000000000) 
    12'h788 : LOC <=          63'b000000000001000000000001000000000000000000000000000000000000000; // D (0x0008008000000000) 
    12'hf13 : LOC <=          63'b000000000001000000000010000000000000000000000000000000000000000; // D (0x0008010000000000) 
    12'hb1c : LOC <=          63'b000000000001000000000100000000000000000000000000000000000000000; // D (0x0008020000000000) 
    12'h302 : LOC <=          63'b000000000001000000001000000000000000000000000000000000000000000; // D (0x0008040000000000) 
    12'h607 : LOC <=          63'b000000000001000000010000000000000000000000000000000000000000000; // D (0x0008080000000000) 
    12'hc0d : LOC <=          63'b000000000001000000100000000000000000000000000000000000000000000; // D (0x0008100000000000) 
    12'hd20 : LOC <=          63'b000000000001000001000000000000000000000000000000000000000000000; // D (0x0008200000000000) 
    12'hf7a : LOC <=          63'b000000000001000010000000000000000000000000000000000000000000000; // D (0x0008400000000000) 
    12'hbce : LOC <=          63'b000000000001000100000000000000000000000000000000000000000000000; // D (0x0008800000000000) 
    12'h2a6 : LOC <=          63'b000000000001001000000000000000000000000000000000000000000000000; // D (0x0009000000000000) 
    12'h54f : LOC <=          63'b000000000001010000000000000000000000000000000000000000000000000; // D (0x000a000000000000) 
    12'ha9d : LOC <=          63'b000000000001100000000000000000000000000000000000000000000000000; // D (0x000c000000000000) 
    12'h001 : LOC <=          63'b000000000001000000000000000000000000000000000000000000000000000; // S (0x0008000000000000) 
//    12'h003 : LOC <=          63'b000000000011000000000000000000000000000000000000000000000000000; // D (0x0018000000000000) 
//    12'h005 : LOC <=          63'b000000000101000000000000000000000000000000000000000000000000000; // D (0x0028000000000000) 
//    12'h009 : LOC <=          63'b000000001001000000000000000000000000000000000000000000000000000; // D (0x0048000000000000) 
//    12'h011 : LOC <=          63'b000000010001000000000000000000000000000000000000000000000000000; // D (0x0088000000000000) 
//    12'h021 : LOC <=          63'b000000100001000000000000000000000000000000000000000000000000000; // D (0x0108000000000000) 
//    12'h041 : LOC <=          63'b000001000001000000000000000000000000000000000000000000000000000; // D (0x0208000000000000) 
//    12'h081 : LOC <=          63'b000010000001000000000000000000000000000000000000000000000000000; // D (0x0408000000000000) 
//    12'h101 : LOC <=          63'b000100000001000000000000000000000000000000000000000000000000000; // D (0x0808000000000000) 
//    12'h201 : LOC <=          63'b001000000001000000000000000000000000000000000000000000000000000; // D (0x1008000000000000) 
//    12'h401 : LOC <=          63'b010000000001000000000000000000000000000000000000000000000000000; // D (0x2008000000000000) 
//    12'h801 : LOC <=          63'b100000000001000000000000000000000000000000000000000000000000000; // D (0x4008000000000000) 
    12'h53b : LOC <=          63'b000000000010000000000000000000000000000000000000000000000000001; // D (0x0010000000000001) 
    12'ha70 : LOC <=          63'b000000000010000000000000000000000000000000000000000000000000010; // D (0x0010000000000002) 
    12'h1df : LOC <=          63'b000000000010000000000000000000000000000000000000000000000000100; // D (0x0010000000000004) 
    12'h3b8 : LOC <=          63'b000000000010000000000000000000000000000000000000000000000001000; // D (0x0010000000000008) 
    12'h776 : LOC <=          63'b000000000010000000000000000000000000000000000000000000000010000; // D (0x0010000000000010) 
    12'heea : LOC <=          63'b000000000010000000000000000000000000000000000000000000000100000; // D (0x0010000000000020) 
    12'h8eb : LOC <=          63'b000000000010000000000000000000000000000000000000000000001000000; // D (0x0010000000000040) 
    12'h4e9 : LOC <=          63'b000000000010000000000000000000000000000000000000000000010000000; // D (0x0010000000000080) 
    12'h9d4 : LOC <=          63'b000000000010000000000000000000000000000000000000000000100000000; // D (0x0010000000000100) 
    12'h697 : LOC <=          63'b000000000010000000000000000000000000000000000000000001000000000; // D (0x0010000000000200) 
    12'hd28 : LOC <=          63'b000000000010000000000000000000000000000000000000000010000000000; // D (0x0010000000000400) 
    12'hf6f : LOC <=          63'b000000000010000000000000000000000000000000000000000100000000000; // D (0x0010000000000800) 
    12'hbe1 : LOC <=          63'b000000000010000000000000000000000000000000000000001000000000000; // D (0x0010000000001000) 
    12'h2fd : LOC <=          63'b000000000010000000000000000000000000000000000000010000000000000; // D (0x0010000000002000) 
    12'h5fc : LOC <=          63'b000000000010000000000000000000000000000000000000100000000000000; // D (0x0010000000004000) 
    12'hbfe : LOC <=          63'b000000000010000000000000000000000000000000000001000000000000000; // D (0x0010000000008000) 
    12'h2c3 : LOC <=          63'b000000000010000000000000000000000000000000000010000000000000000; // D (0x0010000000010000) 
    12'h580 : LOC <=          63'b000000000010000000000000000000000000000000000100000000000000000; // D (0x0010000000020000) 
    12'hb06 : LOC <=          63'b000000000010000000000000000000000000000000001000000000000000000; // D (0x0010000000040000) 
    12'h333 : LOC <=          63'b000000000010000000000000000000000000000000010000000000000000000; // D (0x0010000000080000) 
    12'h660 : LOC <=          63'b000000000010000000000000000000000000000000100000000000000000000; // D (0x0010000000100000) 
    12'hcc6 : LOC <=          63'b000000000010000000000000000000000000000001000000000000000000000; // D (0x0010000000200000) 
    12'hcb3 : LOC <=          63'b000000000010000000000000000000000000000010000000000000000000000; // D (0x0010000000400000) 
    12'hc59 : LOC <=          63'b000000000010000000000000000000000000000100000000000000000000000; // D (0x0010000000800000) 
    12'hd8d : LOC <=          63'b000000000010000000000000000000000000001000000000000000000000000; // D (0x0010000001000000) 
    12'he25 : LOC <=          63'b000000000010000000000000000000000000010000000000000000000000000; // D (0x0010000002000000) 
    12'h975 : LOC <=          63'b000000000010000000000000000000000000100000000000000000000000000; // D (0x0010000004000000) 
    12'h7d5 : LOC <=          63'b000000000010000000000000000000000001000000000000000000000000000; // D (0x0010000008000000) 
    12'hfac : LOC <=          63'b000000000010000000000000000000000010000000000000000000000000000; // D (0x0010000010000000) 
    12'ha67 : LOC <=          63'b000000000010000000000000000000000100000000000000000000000000000; // D (0x0010000020000000) 
    12'h1f1 : LOC <=          63'b000000000010000000000000000000001000000000000000000000000000000; // D (0x0010000040000000) 
    12'h3e4 : LOC <=          63'b000000000010000000000000000000010000000000000000000000000000000; // D (0x0010000080000000) 
    12'h7ce : LOC <=          63'b000000000010000000000000000000100000000000000000000000000000000; // D (0x0010000100000000) 
    12'hf9a : LOC <=          63'b000000000010000000000000000001000000000000000000000000000000000; // D (0x0010000200000000) 
    12'ha0b : LOC <=          63'b000000000010000000000000000010000000000000000000000000000000000; // D (0x0010000400000000) 
    12'h129 : LOC <=          63'b000000000010000000000000000100000000000000000000000000000000000; // D (0x0010000800000000) 
    12'h254 : LOC <=          63'b000000000010000000000000001000000000000000000000000000000000000; // D (0x0010001000000000) 
    12'h4ae : LOC <=          63'b000000000010000000000000010000000000000000000000000000000000000; // D (0x0010002000000000) 
    12'h95a : LOC <=          63'b000000000010000000000000100000000000000000000000000000000000000; // D (0x0010004000000000) 
    12'h78b : LOC <=          63'b000000000010000000000001000000000000000000000000000000000000000; // D (0x0010008000000000) 
    12'hf10 : LOC <=          63'b000000000010000000000010000000000000000000000000000000000000000; // D (0x0010010000000000) 
    12'hb1f : LOC <=          63'b000000000010000000000100000000000000000000000000000000000000000; // D (0x0010020000000000) 
    12'h301 : LOC <=          63'b000000000010000000001000000000000000000000000000000000000000000; // D (0x0010040000000000) 
    12'h604 : LOC <=          63'b000000000010000000010000000000000000000000000000000000000000000; // D (0x0010080000000000) 
    12'hc0e : LOC <=          63'b000000000010000000100000000000000000000000000000000000000000000; // D (0x0010100000000000) 
    12'hd23 : LOC <=          63'b000000000010000001000000000000000000000000000000000000000000000; // D (0x0010200000000000) 
    12'hf79 : LOC <=          63'b000000000010000010000000000000000000000000000000000000000000000; // D (0x0010400000000000) 
    12'hbcd : LOC <=          63'b000000000010000100000000000000000000000000000000000000000000000; // D (0x0010800000000000) 
    12'h2a5 : LOC <=          63'b000000000010001000000000000000000000000000000000000000000000000; // D (0x0011000000000000) 
    12'h54c : LOC <=          63'b000000000010010000000000000000000000000000000000000000000000000; // D (0x0012000000000000) 
    12'ha9e : LOC <=          63'b000000000010100000000000000000000000000000000000000000000000000; // D (0x0014000000000000) 
    12'h003 : LOC <=          63'b000000000011000000000000000000000000000000000000000000000000000; // D (0x0018000000000000) 
    12'h002 : LOC <=          63'b000000000010000000000000000000000000000000000000000000000000000; // S (0x0010000000000000) 
//    12'h006 : LOC <=          63'b000000000110000000000000000000000000000000000000000000000000000; // D (0x0030000000000000) 
//    12'h00a : LOC <=          63'b000000001010000000000000000000000000000000000000000000000000000; // D (0x0050000000000000) 
//    12'h012 : LOC <=          63'b000000010010000000000000000000000000000000000000000000000000000; // D (0x0090000000000000) 
//    12'h022 : LOC <=          63'b000000100010000000000000000000000000000000000000000000000000000; // D (0x0110000000000000) 
//    12'h042 : LOC <=          63'b000001000010000000000000000000000000000000000000000000000000000; // D (0x0210000000000000) 
//    12'h082 : LOC <=          63'b000010000010000000000000000000000000000000000000000000000000000; // D (0x0410000000000000) 
//    12'h102 : LOC <=          63'b000100000010000000000000000000000000000000000000000000000000000; // D (0x0810000000000000) 
//    12'h202 : LOC <=          63'b001000000010000000000000000000000000000000000000000000000000000; // D (0x1010000000000000) 
//    12'h402 : LOC <=          63'b010000000010000000000000000000000000000000000000000000000000000; // D (0x2010000000000000) 
//    12'h802 : LOC <=          63'b100000000010000000000000000000000000000000000000000000000000000; // D (0x4010000000000000) 
    12'h53d : LOC <=          63'b000000000100000000000000000000000000000000000000000000000000001; // D (0x0020000000000001) 
    12'ha76 : LOC <=          63'b000000000100000000000000000000000000000000000000000000000000010; // D (0x0020000000000002) 
    12'h1d9 : LOC <=          63'b000000000100000000000000000000000000000000000000000000000000100; // D (0x0020000000000004) 
    12'h3be : LOC <=          63'b000000000100000000000000000000000000000000000000000000000001000; // D (0x0020000000000008) 
    12'h770 : LOC <=          63'b000000000100000000000000000000000000000000000000000000000010000; // D (0x0020000000000010) 
    12'heec : LOC <=          63'b000000000100000000000000000000000000000000000000000000000100000; // D (0x0020000000000020) 
    12'h8ed : LOC <=          63'b000000000100000000000000000000000000000000000000000000001000000; // D (0x0020000000000040) 
    12'h4ef : LOC <=          63'b000000000100000000000000000000000000000000000000000000010000000; // D (0x0020000000000080) 
    12'h9d2 : LOC <=          63'b000000000100000000000000000000000000000000000000000000100000000; // D (0x0020000000000100) 
    12'h691 : LOC <=          63'b000000000100000000000000000000000000000000000000000001000000000; // D (0x0020000000000200) 
    12'hd2e : LOC <=          63'b000000000100000000000000000000000000000000000000000010000000000; // D (0x0020000000000400) 
    12'hf69 : LOC <=          63'b000000000100000000000000000000000000000000000000000100000000000; // D (0x0020000000000800) 
    12'hbe7 : LOC <=          63'b000000000100000000000000000000000000000000000000001000000000000; // D (0x0020000000001000) 
    12'h2fb : LOC <=          63'b000000000100000000000000000000000000000000000000010000000000000; // D (0x0020000000002000) 
    12'h5fa : LOC <=          63'b000000000100000000000000000000000000000000000000100000000000000; // D (0x0020000000004000) 
    12'hbf8 : LOC <=          63'b000000000100000000000000000000000000000000000001000000000000000; // D (0x0020000000008000) 
    12'h2c5 : LOC <=          63'b000000000100000000000000000000000000000000000010000000000000000; // D (0x0020000000010000) 
    12'h586 : LOC <=          63'b000000000100000000000000000000000000000000000100000000000000000; // D (0x0020000000020000) 
    12'hb00 : LOC <=          63'b000000000100000000000000000000000000000000001000000000000000000; // D (0x0020000000040000) 
    12'h335 : LOC <=          63'b000000000100000000000000000000000000000000010000000000000000000; // D (0x0020000000080000) 
    12'h666 : LOC <=          63'b000000000100000000000000000000000000000000100000000000000000000; // D (0x0020000000100000) 
    12'hcc0 : LOC <=          63'b000000000100000000000000000000000000000001000000000000000000000; // D (0x0020000000200000) 
    12'hcb5 : LOC <=          63'b000000000100000000000000000000000000000010000000000000000000000; // D (0x0020000000400000) 
    12'hc5f : LOC <=          63'b000000000100000000000000000000000000000100000000000000000000000; // D (0x0020000000800000) 
    12'hd8b : LOC <=          63'b000000000100000000000000000000000000001000000000000000000000000; // D (0x0020000001000000) 
    12'he23 : LOC <=          63'b000000000100000000000000000000000000010000000000000000000000000; // D (0x0020000002000000) 
    12'h973 : LOC <=          63'b000000000100000000000000000000000000100000000000000000000000000; // D (0x0020000004000000) 
    12'h7d3 : LOC <=          63'b000000000100000000000000000000000001000000000000000000000000000; // D (0x0020000008000000) 
    12'hfaa : LOC <=          63'b000000000100000000000000000000000010000000000000000000000000000; // D (0x0020000010000000) 
    12'ha61 : LOC <=          63'b000000000100000000000000000000000100000000000000000000000000000; // D (0x0020000020000000) 
    12'h1f7 : LOC <=          63'b000000000100000000000000000000001000000000000000000000000000000; // D (0x0020000040000000) 
    12'h3e2 : LOC <=          63'b000000000100000000000000000000010000000000000000000000000000000; // D (0x0020000080000000) 
    12'h7c8 : LOC <=          63'b000000000100000000000000000000100000000000000000000000000000000; // D (0x0020000100000000) 
    12'hf9c : LOC <=          63'b000000000100000000000000000001000000000000000000000000000000000; // D (0x0020000200000000) 
    12'ha0d : LOC <=          63'b000000000100000000000000000010000000000000000000000000000000000; // D (0x0020000400000000) 
    12'h12f : LOC <=          63'b000000000100000000000000000100000000000000000000000000000000000; // D (0x0020000800000000) 
    12'h252 : LOC <=          63'b000000000100000000000000001000000000000000000000000000000000000; // D (0x0020001000000000) 
    12'h4a8 : LOC <=          63'b000000000100000000000000010000000000000000000000000000000000000; // D (0x0020002000000000) 
    12'h95c : LOC <=          63'b000000000100000000000000100000000000000000000000000000000000000; // D (0x0020004000000000) 
    12'h78d : LOC <=          63'b000000000100000000000001000000000000000000000000000000000000000; // D (0x0020008000000000) 
    12'hf16 : LOC <=          63'b000000000100000000000010000000000000000000000000000000000000000; // D (0x0020010000000000) 
    12'hb19 : LOC <=          63'b000000000100000000000100000000000000000000000000000000000000000; // D (0x0020020000000000) 
    12'h307 : LOC <=          63'b000000000100000000001000000000000000000000000000000000000000000; // D (0x0020040000000000) 
    12'h602 : LOC <=          63'b000000000100000000010000000000000000000000000000000000000000000; // D (0x0020080000000000) 
    12'hc08 : LOC <=          63'b000000000100000000100000000000000000000000000000000000000000000; // D (0x0020100000000000) 
    12'hd25 : LOC <=          63'b000000000100000001000000000000000000000000000000000000000000000; // D (0x0020200000000000) 
    12'hf7f : LOC <=          63'b000000000100000010000000000000000000000000000000000000000000000; // D (0x0020400000000000) 
    12'hbcb : LOC <=          63'b000000000100000100000000000000000000000000000000000000000000000; // D (0x0020800000000000) 
    12'h2a3 : LOC <=          63'b000000000100001000000000000000000000000000000000000000000000000; // D (0x0021000000000000) 
    12'h54a : LOC <=          63'b000000000100010000000000000000000000000000000000000000000000000; // D (0x0022000000000000) 
    12'ha98 : LOC <=          63'b000000000100100000000000000000000000000000000000000000000000000; // D (0x0024000000000000) 
    12'h005 : LOC <=          63'b000000000101000000000000000000000000000000000000000000000000000; // D (0x0028000000000000) 
    12'h006 : LOC <=          63'b000000000110000000000000000000000000000000000000000000000000000; // D (0x0030000000000000) 
    12'h004 : LOC <=          63'b000000000100000000000000000000000000000000000000000000000000000; // S (0x0020000000000000) 
//    12'h00c : LOC <=          63'b000000001100000000000000000000000000000000000000000000000000000; // D (0x0060000000000000) 
//    12'h014 : LOC <=          63'b000000010100000000000000000000000000000000000000000000000000000; // D (0x00a0000000000000) 
//    12'h024 : LOC <=          63'b000000100100000000000000000000000000000000000000000000000000000; // D (0x0120000000000000) 
//    12'h044 : LOC <=          63'b000001000100000000000000000000000000000000000000000000000000000; // D (0x0220000000000000) 
//    12'h084 : LOC <=          63'b000010000100000000000000000000000000000000000000000000000000000; // D (0x0420000000000000) 
//    12'h104 : LOC <=          63'b000100000100000000000000000000000000000000000000000000000000000; // D (0x0820000000000000) 
//    12'h204 : LOC <=          63'b001000000100000000000000000000000000000000000000000000000000000; // D (0x1020000000000000) 
//    12'h404 : LOC <=          63'b010000000100000000000000000000000000000000000000000000000000000; // D (0x2020000000000000) 
//    12'h804 : LOC <=          63'b100000000100000000000000000000000000000000000000000000000000000; // D (0x4020000000000000) 
    12'h531 : LOC <=          63'b000000001000000000000000000000000000000000000000000000000000001; // D (0x0040000000000001) 
    12'ha7a : LOC <=          63'b000000001000000000000000000000000000000000000000000000000000010; // D (0x0040000000000002) 
    12'h1d5 : LOC <=          63'b000000001000000000000000000000000000000000000000000000000000100; // D (0x0040000000000004) 
    12'h3b2 : LOC <=          63'b000000001000000000000000000000000000000000000000000000000001000; // D (0x0040000000000008) 
    12'h77c : LOC <=          63'b000000001000000000000000000000000000000000000000000000000010000; // D (0x0040000000000010) 
    12'hee0 : LOC <=          63'b000000001000000000000000000000000000000000000000000000000100000; // D (0x0040000000000020) 
    12'h8e1 : LOC <=          63'b000000001000000000000000000000000000000000000000000000001000000; // D (0x0040000000000040) 
    12'h4e3 : LOC <=          63'b000000001000000000000000000000000000000000000000000000010000000; // D (0x0040000000000080) 
    12'h9de : LOC <=          63'b000000001000000000000000000000000000000000000000000000100000000; // D (0x0040000000000100) 
    12'h69d : LOC <=          63'b000000001000000000000000000000000000000000000000000001000000000; // D (0x0040000000000200) 
    12'hd22 : LOC <=          63'b000000001000000000000000000000000000000000000000000010000000000; // D (0x0040000000000400) 
    12'hf65 : LOC <=          63'b000000001000000000000000000000000000000000000000000100000000000; // D (0x0040000000000800) 
    12'hbeb : LOC <=          63'b000000001000000000000000000000000000000000000000001000000000000; // D (0x0040000000001000) 
    12'h2f7 : LOC <=          63'b000000001000000000000000000000000000000000000000010000000000000; // D (0x0040000000002000) 
    12'h5f6 : LOC <=          63'b000000001000000000000000000000000000000000000000100000000000000; // D (0x0040000000004000) 
    12'hbf4 : LOC <=          63'b000000001000000000000000000000000000000000000001000000000000000; // D (0x0040000000008000) 
    12'h2c9 : LOC <=          63'b000000001000000000000000000000000000000000000010000000000000000; // D (0x0040000000010000) 
    12'h58a : LOC <=          63'b000000001000000000000000000000000000000000000100000000000000000; // D (0x0040000000020000) 
    12'hb0c : LOC <=          63'b000000001000000000000000000000000000000000001000000000000000000; // D (0x0040000000040000) 
    12'h339 : LOC <=          63'b000000001000000000000000000000000000000000010000000000000000000; // D (0x0040000000080000) 
    12'h66a : LOC <=          63'b000000001000000000000000000000000000000000100000000000000000000; // D (0x0040000000100000) 
    12'hccc : LOC <=          63'b000000001000000000000000000000000000000001000000000000000000000; // D (0x0040000000200000) 
    12'hcb9 : LOC <=          63'b000000001000000000000000000000000000000010000000000000000000000; // D (0x0040000000400000) 
    12'hc53 : LOC <=          63'b000000001000000000000000000000000000000100000000000000000000000; // D (0x0040000000800000) 
    12'hd87 : LOC <=          63'b000000001000000000000000000000000000001000000000000000000000000; // D (0x0040000001000000) 
    12'he2f : LOC <=          63'b000000001000000000000000000000000000010000000000000000000000000; // D (0x0040000002000000) 
    12'h97f : LOC <=          63'b000000001000000000000000000000000000100000000000000000000000000; // D (0x0040000004000000) 
    12'h7df : LOC <=          63'b000000001000000000000000000000000001000000000000000000000000000; // D (0x0040000008000000) 
    12'hfa6 : LOC <=          63'b000000001000000000000000000000000010000000000000000000000000000; // D (0x0040000010000000) 
    12'ha6d : LOC <=          63'b000000001000000000000000000000000100000000000000000000000000000; // D (0x0040000020000000) 
    12'h1fb : LOC <=          63'b000000001000000000000000000000001000000000000000000000000000000; // D (0x0040000040000000) 
    12'h3ee : LOC <=          63'b000000001000000000000000000000010000000000000000000000000000000; // D (0x0040000080000000) 
    12'h7c4 : LOC <=          63'b000000001000000000000000000000100000000000000000000000000000000; // D (0x0040000100000000) 
    12'hf90 : LOC <=          63'b000000001000000000000000000001000000000000000000000000000000000; // D (0x0040000200000000) 
    12'ha01 : LOC <=          63'b000000001000000000000000000010000000000000000000000000000000000; // D (0x0040000400000000) 
    12'h123 : LOC <=          63'b000000001000000000000000000100000000000000000000000000000000000; // D (0x0040000800000000) 
    12'h25e : LOC <=          63'b000000001000000000000000001000000000000000000000000000000000000; // D (0x0040001000000000) 
    12'h4a4 : LOC <=          63'b000000001000000000000000010000000000000000000000000000000000000; // D (0x0040002000000000) 
    12'h950 : LOC <=          63'b000000001000000000000000100000000000000000000000000000000000000; // D (0x0040004000000000) 
    12'h781 : LOC <=          63'b000000001000000000000001000000000000000000000000000000000000000; // D (0x0040008000000000) 
    12'hf1a : LOC <=          63'b000000001000000000000010000000000000000000000000000000000000000; // D (0x0040010000000000) 
    12'hb15 : LOC <=          63'b000000001000000000000100000000000000000000000000000000000000000; // D (0x0040020000000000) 
    12'h30b : LOC <=          63'b000000001000000000001000000000000000000000000000000000000000000; // D (0x0040040000000000) 
    12'h60e : LOC <=          63'b000000001000000000010000000000000000000000000000000000000000000; // D (0x0040080000000000) 
    12'hc04 : LOC <=          63'b000000001000000000100000000000000000000000000000000000000000000; // D (0x0040100000000000) 
    12'hd29 : LOC <=          63'b000000001000000001000000000000000000000000000000000000000000000; // D (0x0040200000000000) 
    12'hf73 : LOC <=          63'b000000001000000010000000000000000000000000000000000000000000000; // D (0x0040400000000000) 
    12'hbc7 : LOC <=          63'b000000001000000100000000000000000000000000000000000000000000000; // D (0x0040800000000000) 
    12'h2af : LOC <=          63'b000000001000001000000000000000000000000000000000000000000000000; // D (0x0041000000000000) 
    12'h546 : LOC <=          63'b000000001000010000000000000000000000000000000000000000000000000; // D (0x0042000000000000) 
    12'ha94 : LOC <=          63'b000000001000100000000000000000000000000000000000000000000000000; // D (0x0044000000000000) 
    12'h009 : LOC <=          63'b000000001001000000000000000000000000000000000000000000000000000; // D (0x0048000000000000) 
    12'h00a : LOC <=          63'b000000001010000000000000000000000000000000000000000000000000000; // D (0x0050000000000000) 
    12'h00c : LOC <=          63'b000000001100000000000000000000000000000000000000000000000000000; // D (0x0060000000000000) 
    12'h008 : LOC <=          63'b000000001000000000000000000000000000000000000000000000000000000; // S (0x0040000000000000) 
//    12'h018 : LOC <=          63'b000000011000000000000000000000000000000000000000000000000000000; // D (0x00c0000000000000) 
//    12'h028 : LOC <=          63'b000000101000000000000000000000000000000000000000000000000000000; // D (0x0140000000000000) 
//    12'h048 : LOC <=          63'b000001001000000000000000000000000000000000000000000000000000000; // D (0x0240000000000000) 
//    12'h088 : LOC <=          63'b000010001000000000000000000000000000000000000000000000000000000; // D (0x0440000000000000) 
//    12'h108 : LOC <=          63'b000100001000000000000000000000000000000000000000000000000000000; // D (0x0840000000000000) 
//    12'h208 : LOC <=          63'b001000001000000000000000000000000000000000000000000000000000000; // D (0x1040000000000000) 
//    12'h408 : LOC <=          63'b010000001000000000000000000000000000000000000000000000000000000; // D (0x2040000000000000) 
//    12'h808 : LOC <=          63'b100000001000000000000000000000000000000000000000000000000000000; // D (0x4040000000000000) 
    12'h529 : LOC <=          63'b000000010000000000000000000000000000000000000000000000000000001; // D (0x0080000000000001) 
    12'ha62 : LOC <=          63'b000000010000000000000000000000000000000000000000000000000000010; // D (0x0080000000000002) 
    12'h1cd : LOC <=          63'b000000010000000000000000000000000000000000000000000000000000100; // D (0x0080000000000004) 
    12'h3aa : LOC <=          63'b000000010000000000000000000000000000000000000000000000000001000; // D (0x0080000000000008) 
    12'h764 : LOC <=          63'b000000010000000000000000000000000000000000000000000000000010000; // D (0x0080000000000010) 
    12'hef8 : LOC <=          63'b000000010000000000000000000000000000000000000000000000000100000; // D (0x0080000000000020) 
    12'h8f9 : LOC <=          63'b000000010000000000000000000000000000000000000000000000001000000; // D (0x0080000000000040) 
    12'h4fb : LOC <=          63'b000000010000000000000000000000000000000000000000000000010000000; // D (0x0080000000000080) 
    12'h9c6 : LOC <=          63'b000000010000000000000000000000000000000000000000000000100000000; // D (0x0080000000000100) 
    12'h685 : LOC <=          63'b000000010000000000000000000000000000000000000000000001000000000; // D (0x0080000000000200) 
    12'hd3a : LOC <=          63'b000000010000000000000000000000000000000000000000000010000000000; // D (0x0080000000000400) 
    12'hf7d : LOC <=          63'b000000010000000000000000000000000000000000000000000100000000000; // D (0x0080000000000800) 
    12'hbf3 : LOC <=          63'b000000010000000000000000000000000000000000000000001000000000000; // D (0x0080000000001000) 
    12'h2ef : LOC <=          63'b000000010000000000000000000000000000000000000000010000000000000; // D (0x0080000000002000) 
    12'h5ee : LOC <=          63'b000000010000000000000000000000000000000000000000100000000000000; // D (0x0080000000004000) 
    12'hbec : LOC <=          63'b000000010000000000000000000000000000000000000001000000000000000; // D (0x0080000000008000) 
    12'h2d1 : LOC <=          63'b000000010000000000000000000000000000000000000010000000000000000; // D (0x0080000000010000) 
    12'h592 : LOC <=          63'b000000010000000000000000000000000000000000000100000000000000000; // D (0x0080000000020000) 
    12'hb14 : LOC <=          63'b000000010000000000000000000000000000000000001000000000000000000; // D (0x0080000000040000) 
    12'h321 : LOC <=          63'b000000010000000000000000000000000000000000010000000000000000000; // D (0x0080000000080000) 
    12'h672 : LOC <=          63'b000000010000000000000000000000000000000000100000000000000000000; // D (0x0080000000100000) 
    12'hcd4 : LOC <=          63'b000000010000000000000000000000000000000001000000000000000000000; // D (0x0080000000200000) 
    12'hca1 : LOC <=          63'b000000010000000000000000000000000000000010000000000000000000000; // D (0x0080000000400000) 
    12'hc4b : LOC <=          63'b000000010000000000000000000000000000000100000000000000000000000; // D (0x0080000000800000) 
    12'hd9f : LOC <=          63'b000000010000000000000000000000000000001000000000000000000000000; // D (0x0080000001000000) 
    12'he37 : LOC <=          63'b000000010000000000000000000000000000010000000000000000000000000; // D (0x0080000002000000) 
    12'h967 : LOC <=          63'b000000010000000000000000000000000000100000000000000000000000000; // D (0x0080000004000000) 
    12'h7c7 : LOC <=          63'b000000010000000000000000000000000001000000000000000000000000000; // D (0x0080000008000000) 
    12'hfbe : LOC <=          63'b000000010000000000000000000000000010000000000000000000000000000; // D (0x0080000010000000) 
    12'ha75 : LOC <=          63'b000000010000000000000000000000000100000000000000000000000000000; // D (0x0080000020000000) 
    12'h1e3 : LOC <=          63'b000000010000000000000000000000001000000000000000000000000000000; // D (0x0080000040000000) 
    12'h3f6 : LOC <=          63'b000000010000000000000000000000010000000000000000000000000000000; // D (0x0080000080000000) 
    12'h7dc : LOC <=          63'b000000010000000000000000000000100000000000000000000000000000000; // D (0x0080000100000000) 
    12'hf88 : LOC <=          63'b000000010000000000000000000001000000000000000000000000000000000; // D (0x0080000200000000) 
    12'ha19 : LOC <=          63'b000000010000000000000000000010000000000000000000000000000000000; // D (0x0080000400000000) 
    12'h13b : LOC <=          63'b000000010000000000000000000100000000000000000000000000000000000; // D (0x0080000800000000) 
    12'h246 : LOC <=          63'b000000010000000000000000001000000000000000000000000000000000000; // D (0x0080001000000000) 
    12'h4bc : LOC <=          63'b000000010000000000000000010000000000000000000000000000000000000; // D (0x0080002000000000) 
    12'h948 : LOC <=          63'b000000010000000000000000100000000000000000000000000000000000000; // D (0x0080004000000000) 
    12'h799 : LOC <=          63'b000000010000000000000001000000000000000000000000000000000000000; // D (0x0080008000000000) 
    12'hf02 : LOC <=          63'b000000010000000000000010000000000000000000000000000000000000000; // D (0x0080010000000000) 
    12'hb0d : LOC <=          63'b000000010000000000000100000000000000000000000000000000000000000; // D (0x0080020000000000) 
    12'h313 : LOC <=          63'b000000010000000000001000000000000000000000000000000000000000000; // D (0x0080040000000000) 
    12'h616 : LOC <=          63'b000000010000000000010000000000000000000000000000000000000000000; // D (0x0080080000000000) 
    12'hc1c : LOC <=          63'b000000010000000000100000000000000000000000000000000000000000000; // D (0x0080100000000000) 
    12'hd31 : LOC <=          63'b000000010000000001000000000000000000000000000000000000000000000; // D (0x0080200000000000) 
    12'hf6b : LOC <=          63'b000000010000000010000000000000000000000000000000000000000000000; // D (0x0080400000000000) 
    12'hbdf : LOC <=          63'b000000010000000100000000000000000000000000000000000000000000000; // D (0x0080800000000000) 
    12'h2b7 : LOC <=          63'b000000010000001000000000000000000000000000000000000000000000000; // D (0x0081000000000000) 
    12'h55e : LOC <=          63'b000000010000010000000000000000000000000000000000000000000000000; // D (0x0082000000000000) 
    12'ha8c : LOC <=          63'b000000010000100000000000000000000000000000000000000000000000000; // D (0x0084000000000000) 
    12'h011 : LOC <=          63'b000000010001000000000000000000000000000000000000000000000000000; // D (0x0088000000000000) 
    12'h012 : LOC <=          63'b000000010010000000000000000000000000000000000000000000000000000; // D (0x0090000000000000) 
    12'h014 : LOC <=          63'b000000010100000000000000000000000000000000000000000000000000000; // D (0x00a0000000000000) 
    12'h018 : LOC <=          63'b000000011000000000000000000000000000000000000000000000000000000; // D (0x00c0000000000000) 
    12'h010 : LOC <=          63'b000000010000000000000000000000000000000000000000000000000000000; // S (0x0080000000000000) 
//    12'h030 : LOC <=          63'b000000110000000000000000000000000000000000000000000000000000000; // D (0x0180000000000000) 
//    12'h050 : LOC <=          63'b000001010000000000000000000000000000000000000000000000000000000; // D (0x0280000000000000) 
//    12'h090 : LOC <=          63'b000010010000000000000000000000000000000000000000000000000000000; // D (0x0480000000000000) 
//    12'h110 : LOC <=          63'b000100010000000000000000000000000000000000000000000000000000000; // D (0x0880000000000000) 
//    12'h210 : LOC <=          63'b001000010000000000000000000000000000000000000000000000000000000; // D (0x1080000000000000) 
//    12'h410 : LOC <=          63'b010000010000000000000000000000000000000000000000000000000000000; // D (0x2080000000000000) 
//    12'h810 : LOC <=          63'b100000010000000000000000000000000000000000000000000000000000000; // D (0x4080000000000000) 
    12'h519 : LOC <=          63'b000000100000000000000000000000000000000000000000000000000000001; // D (0x0100000000000001) 
    12'ha52 : LOC <=          63'b000000100000000000000000000000000000000000000000000000000000010; // D (0x0100000000000002) 
    12'h1fd : LOC <=          63'b000000100000000000000000000000000000000000000000000000000000100; // D (0x0100000000000004) 
    12'h39a : LOC <=          63'b000000100000000000000000000000000000000000000000000000000001000; // D (0x0100000000000008) 
    12'h754 : LOC <=          63'b000000100000000000000000000000000000000000000000000000000010000; // D (0x0100000000000010) 
    12'hec8 : LOC <=          63'b000000100000000000000000000000000000000000000000000000000100000; // D (0x0100000000000020) 
    12'h8c9 : LOC <=          63'b000000100000000000000000000000000000000000000000000000001000000; // D (0x0100000000000040) 
    12'h4cb : LOC <=          63'b000000100000000000000000000000000000000000000000000000010000000; // D (0x0100000000000080) 
    12'h9f6 : LOC <=          63'b000000100000000000000000000000000000000000000000000000100000000; // D (0x0100000000000100) 
    12'h6b5 : LOC <=          63'b000000100000000000000000000000000000000000000000000001000000000; // D (0x0100000000000200) 
    12'hd0a : LOC <=          63'b000000100000000000000000000000000000000000000000000010000000000; // D (0x0100000000000400) 
    12'hf4d : LOC <=          63'b000000100000000000000000000000000000000000000000000100000000000; // D (0x0100000000000800) 
    12'hbc3 : LOC <=          63'b000000100000000000000000000000000000000000000000001000000000000; // D (0x0100000000001000) 
    12'h2df : LOC <=          63'b000000100000000000000000000000000000000000000000010000000000000; // D (0x0100000000002000) 
    12'h5de : LOC <=          63'b000000100000000000000000000000000000000000000000100000000000000; // D (0x0100000000004000) 
    12'hbdc : LOC <=          63'b000000100000000000000000000000000000000000000001000000000000000; // D (0x0100000000008000) 
    12'h2e1 : LOC <=          63'b000000100000000000000000000000000000000000000010000000000000000; // D (0x0100000000010000) 
    12'h5a2 : LOC <=          63'b000000100000000000000000000000000000000000000100000000000000000; // D (0x0100000000020000) 
    12'hb24 : LOC <=          63'b000000100000000000000000000000000000000000001000000000000000000; // D (0x0100000000040000) 
    12'h311 : LOC <=          63'b000000100000000000000000000000000000000000010000000000000000000; // D (0x0100000000080000) 
    12'h642 : LOC <=          63'b000000100000000000000000000000000000000000100000000000000000000; // D (0x0100000000100000) 
    12'hce4 : LOC <=          63'b000000100000000000000000000000000000000001000000000000000000000; // D (0x0100000000200000) 
    12'hc91 : LOC <=          63'b000000100000000000000000000000000000000010000000000000000000000; // D (0x0100000000400000) 
    12'hc7b : LOC <=          63'b000000100000000000000000000000000000000100000000000000000000000; // D (0x0100000000800000) 
    12'hdaf : LOC <=          63'b000000100000000000000000000000000000001000000000000000000000000; // D (0x0100000001000000) 
    12'he07 : LOC <=          63'b000000100000000000000000000000000000010000000000000000000000000; // D (0x0100000002000000) 
    12'h957 : LOC <=          63'b000000100000000000000000000000000000100000000000000000000000000; // D (0x0100000004000000) 
    12'h7f7 : LOC <=          63'b000000100000000000000000000000000001000000000000000000000000000; // D (0x0100000008000000) 
    12'hf8e : LOC <=          63'b000000100000000000000000000000000010000000000000000000000000000; // D (0x0100000010000000) 
    12'ha45 : LOC <=          63'b000000100000000000000000000000000100000000000000000000000000000; // D (0x0100000020000000) 
    12'h1d3 : LOC <=          63'b000000100000000000000000000000001000000000000000000000000000000; // D (0x0100000040000000) 
    12'h3c6 : LOC <=          63'b000000100000000000000000000000010000000000000000000000000000000; // D (0x0100000080000000) 
    12'h7ec : LOC <=          63'b000000100000000000000000000000100000000000000000000000000000000; // D (0x0100000100000000) 
    12'hfb8 : LOC <=          63'b000000100000000000000000000001000000000000000000000000000000000; // D (0x0100000200000000) 
    12'ha29 : LOC <=          63'b000000100000000000000000000010000000000000000000000000000000000; // D (0x0100000400000000) 
    12'h10b : LOC <=          63'b000000100000000000000000000100000000000000000000000000000000000; // D (0x0100000800000000) 
    12'h276 : LOC <=          63'b000000100000000000000000001000000000000000000000000000000000000; // D (0x0100001000000000) 
    12'h48c : LOC <=          63'b000000100000000000000000010000000000000000000000000000000000000; // D (0x0100002000000000) 
    12'h978 : LOC <=          63'b000000100000000000000000100000000000000000000000000000000000000; // D (0x0100004000000000) 
    12'h7a9 : LOC <=          63'b000000100000000000000001000000000000000000000000000000000000000; // D (0x0100008000000000) 
    12'hf32 : LOC <=          63'b000000100000000000000010000000000000000000000000000000000000000; // D (0x0100010000000000) 
    12'hb3d : LOC <=          63'b000000100000000000000100000000000000000000000000000000000000000; // D (0x0100020000000000) 
    12'h323 : LOC <=          63'b000000100000000000001000000000000000000000000000000000000000000; // D (0x0100040000000000) 
    12'h626 : LOC <=          63'b000000100000000000010000000000000000000000000000000000000000000; // D (0x0100080000000000) 
    12'hc2c : LOC <=          63'b000000100000000000100000000000000000000000000000000000000000000; // D (0x0100100000000000) 
    12'hd01 : LOC <=          63'b000000100000000001000000000000000000000000000000000000000000000; // D (0x0100200000000000) 
    12'hf5b : LOC <=          63'b000000100000000010000000000000000000000000000000000000000000000; // D (0x0100400000000000) 
    12'hbef : LOC <=          63'b000000100000000100000000000000000000000000000000000000000000000; // D (0x0100800000000000) 
    12'h287 : LOC <=          63'b000000100000001000000000000000000000000000000000000000000000000; // D (0x0101000000000000) 
    12'h56e : LOC <=          63'b000000100000010000000000000000000000000000000000000000000000000; // D (0x0102000000000000) 
    12'habc : LOC <=          63'b000000100000100000000000000000000000000000000000000000000000000; // D (0x0104000000000000) 
    12'h021 : LOC <=          63'b000000100001000000000000000000000000000000000000000000000000000; // D (0x0108000000000000) 
    12'h022 : LOC <=          63'b000000100010000000000000000000000000000000000000000000000000000; // D (0x0110000000000000) 
    12'h024 : LOC <=          63'b000000100100000000000000000000000000000000000000000000000000000; // D (0x0120000000000000) 
    12'h028 : LOC <=          63'b000000101000000000000000000000000000000000000000000000000000000; // D (0x0140000000000000) 
    12'h030 : LOC <=          63'b000000110000000000000000000000000000000000000000000000000000000; // D (0x0180000000000000) 
    12'h020 : LOC <=          63'b000000100000000000000000000000000000000000000000000000000000000; // S (0x0100000000000000) 
//    12'h060 : LOC <=          63'b000001100000000000000000000000000000000000000000000000000000000; // D (0x0300000000000000) 
//    12'h0a0 : LOC <=          63'b000010100000000000000000000000000000000000000000000000000000000; // D (0x0500000000000000) 
//    12'h120 : LOC <=          63'b000100100000000000000000000000000000000000000000000000000000000; // D (0x0900000000000000) 
//    12'h220 : LOC <=          63'b001000100000000000000000000000000000000000000000000000000000000; // D (0x1100000000000000) 
//    12'h420 : LOC <=          63'b010000100000000000000000000000000000000000000000000000000000000; // D (0x2100000000000000) 
//    12'h820 : LOC <=          63'b100000100000000000000000000000000000000000000000000000000000000; // D (0x4100000000000000) 
    12'h579 : LOC <=          63'b000001000000000000000000000000000000000000000000000000000000001; // D (0x0200000000000001) 
    12'ha32 : LOC <=          63'b000001000000000000000000000000000000000000000000000000000000010; // D (0x0200000000000002) 
    12'h19d : LOC <=          63'b000001000000000000000000000000000000000000000000000000000000100; // D (0x0200000000000004) 
    12'h3fa : LOC <=          63'b000001000000000000000000000000000000000000000000000000000001000; // D (0x0200000000000008) 
    12'h734 : LOC <=          63'b000001000000000000000000000000000000000000000000000000000010000; // D (0x0200000000000010) 
    12'hea8 : LOC <=          63'b000001000000000000000000000000000000000000000000000000000100000; // D (0x0200000000000020) 
    12'h8a9 : LOC <=          63'b000001000000000000000000000000000000000000000000000000001000000; // D (0x0200000000000040) 
    12'h4ab : LOC <=          63'b000001000000000000000000000000000000000000000000000000010000000; // D (0x0200000000000080) 
    12'h996 : LOC <=          63'b000001000000000000000000000000000000000000000000000000100000000; // D (0x0200000000000100) 
    12'h6d5 : LOC <=          63'b000001000000000000000000000000000000000000000000000001000000000; // D (0x0200000000000200) 
    12'hd6a : LOC <=          63'b000001000000000000000000000000000000000000000000000010000000000; // D (0x0200000000000400) 
    12'hf2d : LOC <=          63'b000001000000000000000000000000000000000000000000000100000000000; // D (0x0200000000000800) 
    12'hba3 : LOC <=          63'b000001000000000000000000000000000000000000000000001000000000000; // D (0x0200000000001000) 
    12'h2bf : LOC <=          63'b000001000000000000000000000000000000000000000000010000000000000; // D (0x0200000000002000) 
    12'h5be : LOC <=          63'b000001000000000000000000000000000000000000000000100000000000000; // D (0x0200000000004000) 
    12'hbbc : LOC <=          63'b000001000000000000000000000000000000000000000001000000000000000; // D (0x0200000000008000) 
    12'h281 : LOC <=          63'b000001000000000000000000000000000000000000000010000000000000000; // D (0x0200000000010000) 
    12'h5c2 : LOC <=          63'b000001000000000000000000000000000000000000000100000000000000000; // D (0x0200000000020000) 
    12'hb44 : LOC <=          63'b000001000000000000000000000000000000000000001000000000000000000; // D (0x0200000000040000) 
    12'h371 : LOC <=          63'b000001000000000000000000000000000000000000010000000000000000000; // D (0x0200000000080000) 
    12'h622 : LOC <=          63'b000001000000000000000000000000000000000000100000000000000000000; // D (0x0200000000100000) 
    12'hc84 : LOC <=          63'b000001000000000000000000000000000000000001000000000000000000000; // D (0x0200000000200000) 
    12'hcf1 : LOC <=          63'b000001000000000000000000000000000000000010000000000000000000000; // D (0x0200000000400000) 
    12'hc1b : LOC <=          63'b000001000000000000000000000000000000000100000000000000000000000; // D (0x0200000000800000) 
    12'hdcf : LOC <=          63'b000001000000000000000000000000000000001000000000000000000000000; // D (0x0200000001000000) 
    12'he67 : LOC <=          63'b000001000000000000000000000000000000010000000000000000000000000; // D (0x0200000002000000) 
    12'h937 : LOC <=          63'b000001000000000000000000000000000000100000000000000000000000000; // D (0x0200000004000000) 
    12'h797 : LOC <=          63'b000001000000000000000000000000000001000000000000000000000000000; // D (0x0200000008000000) 
    12'hfee : LOC <=          63'b000001000000000000000000000000000010000000000000000000000000000; // D (0x0200000010000000) 
    12'ha25 : LOC <=          63'b000001000000000000000000000000000100000000000000000000000000000; // D (0x0200000020000000) 
    12'h1b3 : LOC <=          63'b000001000000000000000000000000001000000000000000000000000000000; // D (0x0200000040000000) 
    12'h3a6 : LOC <=          63'b000001000000000000000000000000010000000000000000000000000000000; // D (0x0200000080000000) 
    12'h78c : LOC <=          63'b000001000000000000000000000000100000000000000000000000000000000; // D (0x0200000100000000) 
    12'hfd8 : LOC <=          63'b000001000000000000000000000001000000000000000000000000000000000; // D (0x0200000200000000) 
    12'ha49 : LOC <=          63'b000001000000000000000000000010000000000000000000000000000000000; // D (0x0200000400000000) 
    12'h16b : LOC <=          63'b000001000000000000000000000100000000000000000000000000000000000; // D (0x0200000800000000) 
    12'h216 : LOC <=          63'b000001000000000000000000001000000000000000000000000000000000000; // D (0x0200001000000000) 
    12'h4ec : LOC <=          63'b000001000000000000000000010000000000000000000000000000000000000; // D (0x0200002000000000) 
    12'h918 : LOC <=          63'b000001000000000000000000100000000000000000000000000000000000000; // D (0x0200004000000000) 
    12'h7c9 : LOC <=          63'b000001000000000000000001000000000000000000000000000000000000000; // D (0x0200008000000000) 
    12'hf52 : LOC <=          63'b000001000000000000000010000000000000000000000000000000000000000; // D (0x0200010000000000) 
    12'hb5d : LOC <=          63'b000001000000000000000100000000000000000000000000000000000000000; // D (0x0200020000000000) 
    12'h343 : LOC <=          63'b000001000000000000001000000000000000000000000000000000000000000; // D (0x0200040000000000) 
    12'h646 : LOC <=          63'b000001000000000000010000000000000000000000000000000000000000000; // D (0x0200080000000000) 
    12'hc4c : LOC <=          63'b000001000000000000100000000000000000000000000000000000000000000; // D (0x0200100000000000) 
    12'hd61 : LOC <=          63'b000001000000000001000000000000000000000000000000000000000000000; // D (0x0200200000000000) 
    12'hf3b : LOC <=          63'b000001000000000010000000000000000000000000000000000000000000000; // D (0x0200400000000000) 
    12'hb8f : LOC <=          63'b000001000000000100000000000000000000000000000000000000000000000; // D (0x0200800000000000) 
    12'h2e7 : LOC <=          63'b000001000000001000000000000000000000000000000000000000000000000; // D (0x0201000000000000) 
    12'h50e : LOC <=          63'b000001000000010000000000000000000000000000000000000000000000000; // D (0x0202000000000000) 
    12'hadc : LOC <=          63'b000001000000100000000000000000000000000000000000000000000000000; // D (0x0204000000000000) 
    12'h041 : LOC <=          63'b000001000001000000000000000000000000000000000000000000000000000; // D (0x0208000000000000) 
    12'h042 : LOC <=          63'b000001000010000000000000000000000000000000000000000000000000000; // D (0x0210000000000000) 
    12'h044 : LOC <=          63'b000001000100000000000000000000000000000000000000000000000000000; // D (0x0220000000000000) 
    12'h048 : LOC <=          63'b000001001000000000000000000000000000000000000000000000000000000; // D (0x0240000000000000) 
    12'h050 : LOC <=          63'b000001010000000000000000000000000000000000000000000000000000000; // D (0x0280000000000000) 
    12'h060 : LOC <=          63'b000001100000000000000000000000000000000000000000000000000000000; // D (0x0300000000000000) 
    12'h040 : LOC <=          63'b000001000000000000000000000000000000000000000000000000000000000; // S (0x0200000000000000) 
//    12'h0c0 : LOC <=          63'b000011000000000000000000000000000000000000000000000000000000000; // D (0x0600000000000000) 
//    12'h140 : LOC <=          63'b000101000000000000000000000000000000000000000000000000000000000; // D (0x0a00000000000000) 
//    12'h240 : LOC <=          63'b001001000000000000000000000000000000000000000000000000000000000; // D (0x1200000000000000) 
//    12'h440 : LOC <=          63'b010001000000000000000000000000000000000000000000000000000000000; // D (0x2200000000000000) 
//    12'h840 : LOC <=          63'b100001000000000000000000000000000000000000000000000000000000000; // D (0x4200000000000000) 
    12'h5b9 : LOC <=          63'b000010000000000000000000000000000000000000000000000000000000001; // D (0x0400000000000001) 
    12'haf2 : LOC <=          63'b000010000000000000000000000000000000000000000000000000000000010; // D (0x0400000000000002) 
    12'h15d : LOC <=          63'b000010000000000000000000000000000000000000000000000000000000100; // D (0x0400000000000004) 
    12'h33a : LOC <=          63'b000010000000000000000000000000000000000000000000000000000001000; // D (0x0400000000000008) 
    12'h7f4 : LOC <=          63'b000010000000000000000000000000000000000000000000000000000010000; // D (0x0400000000000010) 
    12'he68 : LOC <=          63'b000010000000000000000000000000000000000000000000000000000100000; // D (0x0400000000000020) 
    12'h869 : LOC <=          63'b000010000000000000000000000000000000000000000000000000001000000; // D (0x0400000000000040) 
    12'h46b : LOC <=          63'b000010000000000000000000000000000000000000000000000000010000000; // D (0x0400000000000080) 
    12'h956 : LOC <=          63'b000010000000000000000000000000000000000000000000000000100000000; // D (0x0400000000000100) 
    12'h615 : LOC <=          63'b000010000000000000000000000000000000000000000000000001000000000; // D (0x0400000000000200) 
    12'hdaa : LOC <=          63'b000010000000000000000000000000000000000000000000000010000000000; // D (0x0400000000000400) 
    12'hfed : LOC <=          63'b000010000000000000000000000000000000000000000000000100000000000; // D (0x0400000000000800) 
    12'hb63 : LOC <=          63'b000010000000000000000000000000000000000000000000001000000000000; // D (0x0400000000001000) 
    12'h27f : LOC <=          63'b000010000000000000000000000000000000000000000000010000000000000; // D (0x0400000000002000) 
    12'h57e : LOC <=          63'b000010000000000000000000000000000000000000000000100000000000000; // D (0x0400000000004000) 
    12'hb7c : LOC <=          63'b000010000000000000000000000000000000000000000001000000000000000; // D (0x0400000000008000) 
    12'h241 : LOC <=          63'b000010000000000000000000000000000000000000000010000000000000000; // D (0x0400000000010000) 
    12'h502 : LOC <=          63'b000010000000000000000000000000000000000000000100000000000000000; // D (0x0400000000020000) 
    12'hb84 : LOC <=          63'b000010000000000000000000000000000000000000001000000000000000000; // D (0x0400000000040000) 
    12'h3b1 : LOC <=          63'b000010000000000000000000000000000000000000010000000000000000000; // D (0x0400000000080000) 
    12'h6e2 : LOC <=          63'b000010000000000000000000000000000000000000100000000000000000000; // D (0x0400000000100000) 
    12'hc44 : LOC <=          63'b000010000000000000000000000000000000000001000000000000000000000; // D (0x0400000000200000) 
    12'hc31 : LOC <=          63'b000010000000000000000000000000000000000010000000000000000000000; // D (0x0400000000400000) 
    12'hcdb : LOC <=          63'b000010000000000000000000000000000000000100000000000000000000000; // D (0x0400000000800000) 
    12'hd0f : LOC <=          63'b000010000000000000000000000000000000001000000000000000000000000; // D (0x0400000001000000) 
    12'hea7 : LOC <=          63'b000010000000000000000000000000000000010000000000000000000000000; // D (0x0400000002000000) 
    12'h9f7 : LOC <=          63'b000010000000000000000000000000000000100000000000000000000000000; // D (0x0400000004000000) 
    12'h757 : LOC <=          63'b000010000000000000000000000000000001000000000000000000000000000; // D (0x0400000008000000) 
    12'hf2e : LOC <=          63'b000010000000000000000000000000000010000000000000000000000000000; // D (0x0400000010000000) 
    12'hae5 : LOC <=          63'b000010000000000000000000000000000100000000000000000000000000000; // D (0x0400000020000000) 
    12'h173 : LOC <=          63'b000010000000000000000000000000001000000000000000000000000000000; // D (0x0400000040000000) 
    12'h366 : LOC <=          63'b000010000000000000000000000000010000000000000000000000000000000; // D (0x0400000080000000) 
    12'h74c : LOC <=          63'b000010000000000000000000000000100000000000000000000000000000000; // D (0x0400000100000000) 
    12'hf18 : LOC <=          63'b000010000000000000000000000001000000000000000000000000000000000; // D (0x0400000200000000) 
    12'ha89 : LOC <=          63'b000010000000000000000000000010000000000000000000000000000000000; // D (0x0400000400000000) 
    12'h1ab : LOC <=          63'b000010000000000000000000000100000000000000000000000000000000000; // D (0x0400000800000000) 
    12'h2d6 : LOC <=          63'b000010000000000000000000001000000000000000000000000000000000000; // D (0x0400001000000000) 
    12'h42c : LOC <=          63'b000010000000000000000000010000000000000000000000000000000000000; // D (0x0400002000000000) 
    12'h9d8 : LOC <=          63'b000010000000000000000000100000000000000000000000000000000000000; // D (0x0400004000000000) 
    12'h709 : LOC <=          63'b000010000000000000000001000000000000000000000000000000000000000; // D (0x0400008000000000) 
    12'hf92 : LOC <=          63'b000010000000000000000010000000000000000000000000000000000000000; // D (0x0400010000000000) 
    12'hb9d : LOC <=          63'b000010000000000000000100000000000000000000000000000000000000000; // D (0x0400020000000000) 
    12'h383 : LOC <=          63'b000010000000000000001000000000000000000000000000000000000000000; // D (0x0400040000000000) 
    12'h686 : LOC <=          63'b000010000000000000010000000000000000000000000000000000000000000; // D (0x0400080000000000) 
    12'hc8c : LOC <=          63'b000010000000000000100000000000000000000000000000000000000000000; // D (0x0400100000000000) 
    12'hda1 : LOC <=          63'b000010000000000001000000000000000000000000000000000000000000000; // D (0x0400200000000000) 
    12'hffb : LOC <=          63'b000010000000000010000000000000000000000000000000000000000000000; // D (0x0400400000000000) 
    12'hb4f : LOC <=          63'b000010000000000100000000000000000000000000000000000000000000000; // D (0x0400800000000000) 
    12'h227 : LOC <=          63'b000010000000001000000000000000000000000000000000000000000000000; // D (0x0401000000000000) 
    12'h5ce : LOC <=          63'b000010000000010000000000000000000000000000000000000000000000000; // D (0x0402000000000000) 
    12'ha1c : LOC <=          63'b000010000000100000000000000000000000000000000000000000000000000; // D (0x0404000000000000) 
    12'h081 : LOC <=          63'b000010000001000000000000000000000000000000000000000000000000000; // D (0x0408000000000000) 
    12'h082 : LOC <=          63'b000010000010000000000000000000000000000000000000000000000000000; // D (0x0410000000000000) 
    12'h084 : LOC <=          63'b000010000100000000000000000000000000000000000000000000000000000; // D (0x0420000000000000) 
    12'h088 : LOC <=          63'b000010001000000000000000000000000000000000000000000000000000000; // D (0x0440000000000000) 
    12'h090 : LOC <=          63'b000010010000000000000000000000000000000000000000000000000000000; // D (0x0480000000000000) 
    12'h0a0 : LOC <=          63'b000010100000000000000000000000000000000000000000000000000000000; // D (0x0500000000000000) 
    12'h0c0 : LOC <=          63'b000011000000000000000000000000000000000000000000000000000000000; // D (0x0600000000000000) 
    12'h080 : LOC <=          63'b000010000000000000000000000000000000000000000000000000000000000; // S (0x0400000000000000) 
//    12'h180 : LOC <=          63'b000110000000000000000000000000000000000000000000000000000000000; // D (0x0c00000000000000) 
//    12'h280 : LOC <=          63'b001010000000000000000000000000000000000000000000000000000000000; // D (0x1400000000000000) 
//    12'h480 : LOC <=          63'b010010000000000000000000000000000000000000000000000000000000000; // D (0x2400000000000000) 
//    12'h880 : LOC <=          63'b100010000000000000000000000000000000000000000000000000000000000; // D (0x4400000000000000) 
    12'h439 : LOC <=          63'b000100000000000000000000000000000000000000000000000000000000001; // D (0x0800000000000001) 
    12'hb72 : LOC <=          63'b000100000000000000000000000000000000000000000000000000000000010; // D (0x0800000000000002) 
    12'h0dd : LOC <=          63'b000100000000000000000000000000000000000000000000000000000000100; // D (0x0800000000000004) 
    12'h2ba : LOC <=          63'b000100000000000000000000000000000000000000000000000000000001000; // D (0x0800000000000008) 
    12'h674 : LOC <=          63'b000100000000000000000000000000000000000000000000000000000010000; // D (0x0800000000000010) 
    12'hfe8 : LOC <=          63'b000100000000000000000000000000000000000000000000000000000100000; // D (0x0800000000000020) 
    12'h9e9 : LOC <=          63'b000100000000000000000000000000000000000000000000000000001000000; // D (0x0800000000000040) 
    12'h5eb : LOC <=          63'b000100000000000000000000000000000000000000000000000000010000000; // D (0x0800000000000080) 
    12'h8d6 : LOC <=          63'b000100000000000000000000000000000000000000000000000000100000000; // D (0x0800000000000100) 
    12'h795 : LOC <=          63'b000100000000000000000000000000000000000000000000000001000000000; // D (0x0800000000000200) 
    12'hc2a : LOC <=          63'b000100000000000000000000000000000000000000000000000010000000000; // D (0x0800000000000400) 
    12'he6d : LOC <=          63'b000100000000000000000000000000000000000000000000000100000000000; // D (0x0800000000000800) 
    12'hae3 : LOC <=          63'b000100000000000000000000000000000000000000000000001000000000000; // D (0x0800000000001000) 
    12'h3ff : LOC <=          63'b000100000000000000000000000000000000000000000000010000000000000; // D (0x0800000000002000) 
    12'h4fe : LOC <=          63'b000100000000000000000000000000000000000000000000100000000000000; // D (0x0800000000004000) 
    12'hafc : LOC <=          63'b000100000000000000000000000000000000000000000001000000000000000; // D (0x0800000000008000) 
    12'h3c1 : LOC <=          63'b000100000000000000000000000000000000000000000010000000000000000; // D (0x0800000000010000) 
    12'h482 : LOC <=          63'b000100000000000000000000000000000000000000000100000000000000000; // D (0x0800000000020000) 
    12'ha04 : LOC <=          63'b000100000000000000000000000000000000000000001000000000000000000; // D (0x0800000000040000) 
    12'h231 : LOC <=          63'b000100000000000000000000000000000000000000010000000000000000000; // D (0x0800000000080000) 
    12'h762 : LOC <=          63'b000100000000000000000000000000000000000000100000000000000000000; // D (0x0800000000100000) 
    12'hdc4 : LOC <=          63'b000100000000000000000000000000000000000001000000000000000000000; // D (0x0800000000200000) 
    12'hdb1 : LOC <=          63'b000100000000000000000000000000000000000010000000000000000000000; // D (0x0800000000400000) 
    12'hd5b : LOC <=          63'b000100000000000000000000000000000000000100000000000000000000000; // D (0x0800000000800000) 
    12'hc8f : LOC <=          63'b000100000000000000000000000000000000001000000000000000000000000; // D (0x0800000001000000) 
    12'hf27 : LOC <=          63'b000100000000000000000000000000000000010000000000000000000000000; // D (0x0800000002000000) 
    12'h877 : LOC <=          63'b000100000000000000000000000000000000100000000000000000000000000; // D (0x0800000004000000) 
    12'h6d7 : LOC <=          63'b000100000000000000000000000000000001000000000000000000000000000; // D (0x0800000008000000) 
    12'heae : LOC <=          63'b000100000000000000000000000000000010000000000000000000000000000; // D (0x0800000010000000) 
    12'hb65 : LOC <=          63'b000100000000000000000000000000000100000000000000000000000000000; // D (0x0800000020000000) 
    12'h0f3 : LOC <=          63'b000100000000000000000000000000001000000000000000000000000000000; // D (0x0800000040000000) 
    12'h2e6 : LOC <=          63'b000100000000000000000000000000010000000000000000000000000000000; // D (0x0800000080000000) 
    12'h6cc : LOC <=          63'b000100000000000000000000000000100000000000000000000000000000000; // D (0x0800000100000000) 
    12'he98 : LOC <=          63'b000100000000000000000000000001000000000000000000000000000000000; // D (0x0800000200000000) 
    12'hb09 : LOC <=          63'b000100000000000000000000000010000000000000000000000000000000000; // D (0x0800000400000000) 
    12'h02b : LOC <=          63'b000100000000000000000000000100000000000000000000000000000000000; // D (0x0800000800000000) 
    12'h356 : LOC <=          63'b000100000000000000000000001000000000000000000000000000000000000; // D (0x0800001000000000) 
    12'h5ac : LOC <=          63'b000100000000000000000000010000000000000000000000000000000000000; // D (0x0800002000000000) 
    12'h858 : LOC <=          63'b000100000000000000000000100000000000000000000000000000000000000; // D (0x0800004000000000) 
    12'h689 : LOC <=          63'b000100000000000000000001000000000000000000000000000000000000000; // D (0x0800008000000000) 
    12'he12 : LOC <=          63'b000100000000000000000010000000000000000000000000000000000000000; // D (0x0800010000000000) 
    12'ha1d : LOC <=          63'b000100000000000000000100000000000000000000000000000000000000000; // D (0x0800020000000000) 
    12'h203 : LOC <=          63'b000100000000000000001000000000000000000000000000000000000000000; // D (0x0800040000000000) 
    12'h706 : LOC <=          63'b000100000000000000010000000000000000000000000000000000000000000; // D (0x0800080000000000) 
    12'hd0c : LOC <=          63'b000100000000000000100000000000000000000000000000000000000000000; // D (0x0800100000000000) 
    12'hc21 : LOC <=          63'b000100000000000001000000000000000000000000000000000000000000000; // D (0x0800200000000000) 
    12'he7b : LOC <=          63'b000100000000000010000000000000000000000000000000000000000000000; // D (0x0800400000000000) 
    12'hacf : LOC <=          63'b000100000000000100000000000000000000000000000000000000000000000; // D (0x0800800000000000) 
    12'h3a7 : LOC <=          63'b000100000000001000000000000000000000000000000000000000000000000; // D (0x0801000000000000) 
    12'h44e : LOC <=          63'b000100000000010000000000000000000000000000000000000000000000000; // D (0x0802000000000000) 
    12'hb9c : LOC <=          63'b000100000000100000000000000000000000000000000000000000000000000; // D (0x0804000000000000) 
    12'h101 : LOC <=          63'b000100000001000000000000000000000000000000000000000000000000000; // D (0x0808000000000000) 
    12'h102 : LOC <=          63'b000100000010000000000000000000000000000000000000000000000000000; // D (0x0810000000000000) 
    12'h104 : LOC <=          63'b000100000100000000000000000000000000000000000000000000000000000; // D (0x0820000000000000) 
    12'h108 : LOC <=          63'b000100001000000000000000000000000000000000000000000000000000000; // D (0x0840000000000000) 
    12'h110 : LOC <=          63'b000100010000000000000000000000000000000000000000000000000000000; // D (0x0880000000000000) 
    12'h120 : LOC <=          63'b000100100000000000000000000000000000000000000000000000000000000; // D (0x0900000000000000) 
    12'h140 : LOC <=          63'b000101000000000000000000000000000000000000000000000000000000000; // D (0x0a00000000000000) 
    12'h180 : LOC <=          63'b000110000000000000000000000000000000000000000000000000000000000; // D (0x0c00000000000000) 
    12'h100 : LOC <=          63'b000100000000000000000000000000000000000000000000000000000000000; // S (0x0800000000000000) 
//    12'h300 : LOC <=          63'b001100000000000000000000000000000000000000000000000000000000000; // D (0x1800000000000000) 
//    12'h500 : LOC <=          63'b010100000000000000000000000000000000000000000000000000000000000; // D (0x2800000000000000) 
//    12'h900 : LOC <=          63'b100100000000000000000000000000000000000000000000000000000000000; // D (0x4800000000000000) 
    12'h739 : LOC <=          63'b001000000000000000000000000000000000000000000000000000000000001; // D (0x1000000000000001) 
    12'h872 : LOC <=          63'b001000000000000000000000000000000000000000000000000000000000010; // D (0x1000000000000002) 
    12'h3dd : LOC <=          63'b001000000000000000000000000000000000000000000000000000000000100; // D (0x1000000000000004) 
    12'h1ba : LOC <=          63'b001000000000000000000000000000000000000000000000000000000001000; // D (0x1000000000000008) 
    12'h574 : LOC <=          63'b001000000000000000000000000000000000000000000000000000000010000; // D (0x1000000000000010) 
    12'hce8 : LOC <=          63'b001000000000000000000000000000000000000000000000000000000100000; // D (0x1000000000000020) 
    12'hae9 : LOC <=          63'b001000000000000000000000000000000000000000000000000000001000000; // D (0x1000000000000040) 
    12'h6eb : LOC <=          63'b001000000000000000000000000000000000000000000000000000010000000; // D (0x1000000000000080) 
    12'hbd6 : LOC <=          63'b001000000000000000000000000000000000000000000000000000100000000; // D (0x1000000000000100) 
    12'h495 : LOC <=          63'b001000000000000000000000000000000000000000000000000001000000000; // D (0x1000000000000200) 
    12'hf2a : LOC <=          63'b001000000000000000000000000000000000000000000000000010000000000; // D (0x1000000000000400) 
    12'hd6d : LOC <=          63'b001000000000000000000000000000000000000000000000000100000000000; // D (0x1000000000000800) 
    12'h9e3 : LOC <=          63'b001000000000000000000000000000000000000000000000001000000000000; // D (0x1000000000001000) 
    12'h0ff : LOC <=          63'b001000000000000000000000000000000000000000000000010000000000000; // D (0x1000000000002000) 
    12'h7fe : LOC <=          63'b001000000000000000000000000000000000000000000000100000000000000; // D (0x1000000000004000) 
    12'h9fc : LOC <=          63'b001000000000000000000000000000000000000000000001000000000000000; // D (0x1000000000008000) 
    12'h0c1 : LOC <=          63'b001000000000000000000000000000000000000000000010000000000000000; // D (0x1000000000010000) 
    12'h782 : LOC <=          63'b001000000000000000000000000000000000000000000100000000000000000; // D (0x1000000000020000) 
    12'h904 : LOC <=          63'b001000000000000000000000000000000000000000001000000000000000000; // D (0x1000000000040000) 
    12'h131 : LOC <=          63'b001000000000000000000000000000000000000000010000000000000000000; // D (0x1000000000080000) 
    12'h462 : LOC <=          63'b001000000000000000000000000000000000000000100000000000000000000; // D (0x1000000000100000) 
    12'hec4 : LOC <=          63'b001000000000000000000000000000000000000001000000000000000000000; // D (0x1000000000200000) 
    12'heb1 : LOC <=          63'b001000000000000000000000000000000000000010000000000000000000000; // D (0x1000000000400000) 
    12'he5b : LOC <=          63'b001000000000000000000000000000000000000100000000000000000000000; // D (0x1000000000800000) 
    12'hf8f : LOC <=          63'b001000000000000000000000000000000000001000000000000000000000000; // D (0x1000000001000000) 
    12'hc27 : LOC <=          63'b001000000000000000000000000000000000010000000000000000000000000; // D (0x1000000002000000) 
    12'hb77 : LOC <=          63'b001000000000000000000000000000000000100000000000000000000000000; // D (0x1000000004000000) 
    12'h5d7 : LOC <=          63'b001000000000000000000000000000000001000000000000000000000000000; // D (0x1000000008000000) 
    12'hdae : LOC <=          63'b001000000000000000000000000000000010000000000000000000000000000; // D (0x1000000010000000) 
    12'h865 : LOC <=          63'b001000000000000000000000000000000100000000000000000000000000000; // D (0x1000000020000000) 
    12'h3f3 : LOC <=          63'b001000000000000000000000000000001000000000000000000000000000000; // D (0x1000000040000000) 
    12'h1e6 : LOC <=          63'b001000000000000000000000000000010000000000000000000000000000000; // D (0x1000000080000000) 
    12'h5cc : LOC <=          63'b001000000000000000000000000000100000000000000000000000000000000; // D (0x1000000100000000) 
    12'hd98 : LOC <=          63'b001000000000000000000000000001000000000000000000000000000000000; // D (0x1000000200000000) 
    12'h809 : LOC <=          63'b001000000000000000000000000010000000000000000000000000000000000; // D (0x1000000400000000) 
    12'h32b : LOC <=          63'b001000000000000000000000000100000000000000000000000000000000000; // D (0x1000000800000000) 
    12'h056 : LOC <=          63'b001000000000000000000000001000000000000000000000000000000000000; // D (0x1000001000000000) 
    12'h6ac : LOC <=          63'b001000000000000000000000010000000000000000000000000000000000000; // D (0x1000002000000000) 
    12'hb58 : LOC <=          63'b001000000000000000000000100000000000000000000000000000000000000; // D (0x1000004000000000) 
    12'h589 : LOC <=          63'b001000000000000000000001000000000000000000000000000000000000000; // D (0x1000008000000000) 
    12'hd12 : LOC <=          63'b001000000000000000000010000000000000000000000000000000000000000; // D (0x1000010000000000) 
    12'h91d : LOC <=          63'b001000000000000000000100000000000000000000000000000000000000000; // D (0x1000020000000000) 
    12'h103 : LOC <=          63'b001000000000000000001000000000000000000000000000000000000000000; // D (0x1000040000000000) 
    12'h406 : LOC <=          63'b001000000000000000010000000000000000000000000000000000000000000; // D (0x1000080000000000) 
    12'he0c : LOC <=          63'b001000000000000000100000000000000000000000000000000000000000000; // D (0x1000100000000000) 
    12'hf21 : LOC <=          63'b001000000000000001000000000000000000000000000000000000000000000; // D (0x1000200000000000) 
    12'hd7b : LOC <=          63'b001000000000000010000000000000000000000000000000000000000000000; // D (0x1000400000000000) 
    12'h9cf : LOC <=          63'b001000000000000100000000000000000000000000000000000000000000000; // D (0x1000800000000000) 
    12'h0a7 : LOC <=          63'b001000000000001000000000000000000000000000000000000000000000000; // D (0x1001000000000000) 
    12'h74e : LOC <=          63'b001000000000010000000000000000000000000000000000000000000000000; // D (0x1002000000000000) 
    12'h89c : LOC <=          63'b001000000000100000000000000000000000000000000000000000000000000; // D (0x1004000000000000) 
    12'h201 : LOC <=          63'b001000000001000000000000000000000000000000000000000000000000000; // D (0x1008000000000000) 
    12'h202 : LOC <=          63'b001000000010000000000000000000000000000000000000000000000000000; // D (0x1010000000000000) 
    12'h204 : LOC <=          63'b001000000100000000000000000000000000000000000000000000000000000; // D (0x1020000000000000) 
    12'h208 : LOC <=          63'b001000001000000000000000000000000000000000000000000000000000000; // D (0x1040000000000000) 
    12'h210 : LOC <=          63'b001000010000000000000000000000000000000000000000000000000000000; // D (0x1080000000000000) 
    12'h220 : LOC <=          63'b001000100000000000000000000000000000000000000000000000000000000; // D (0x1100000000000000) 
    12'h240 : LOC <=          63'b001001000000000000000000000000000000000000000000000000000000000; // D (0x1200000000000000) 
    12'h280 : LOC <=          63'b001010000000000000000000000000000000000000000000000000000000000; // D (0x1400000000000000) 
    12'h300 : LOC <=          63'b001100000000000000000000000000000000000000000000000000000000000; // D (0x1800000000000000) 
    12'h200 : LOC <=          63'b001000000000000000000000000000000000000000000000000000000000000; // S (0x1000000000000000) 
//    12'h600 : LOC <=          63'b011000000000000000000000000000000000000000000000000000000000000; // D (0x3000000000000000) 
//    12'ha00 : LOC <=          63'b101000000000000000000000000000000000000000000000000000000000000; // D (0x5000000000000000) 
    12'h139 : LOC <=          63'b010000000000000000000000000000000000000000000000000000000000001; // D (0x2000000000000001) 
    12'he72 : LOC <=          63'b010000000000000000000000000000000000000000000000000000000000010; // D (0x2000000000000002) 
    12'h5dd : LOC <=          63'b010000000000000000000000000000000000000000000000000000000000100; // D (0x2000000000000004) 
    12'h7ba : LOC <=          63'b010000000000000000000000000000000000000000000000000000000001000; // D (0x2000000000000008) 
    12'h374 : LOC <=          63'b010000000000000000000000000000000000000000000000000000000010000; // D (0x2000000000000010) 
    12'hae8 : LOC <=          63'b010000000000000000000000000000000000000000000000000000000100000; // D (0x2000000000000020) 
    12'hce9 : LOC <=          63'b010000000000000000000000000000000000000000000000000000001000000; // D (0x2000000000000040) 
    12'h0eb : LOC <=          63'b010000000000000000000000000000000000000000000000000000010000000; // D (0x2000000000000080) 
    12'hdd6 : LOC <=          63'b010000000000000000000000000000000000000000000000000000100000000; // D (0x2000000000000100) 
    12'h295 : LOC <=          63'b010000000000000000000000000000000000000000000000000001000000000; // D (0x2000000000000200) 
    12'h92a : LOC <=          63'b010000000000000000000000000000000000000000000000000010000000000; // D (0x2000000000000400) 
    12'hb6d : LOC <=          63'b010000000000000000000000000000000000000000000000000100000000000; // D (0x2000000000000800) 
    12'hfe3 : LOC <=          63'b010000000000000000000000000000000000000000000000001000000000000; // D (0x2000000000001000) 
    12'h6ff : LOC <=          63'b010000000000000000000000000000000000000000000000010000000000000; // D (0x2000000000002000) 
    12'h1fe : LOC <=          63'b010000000000000000000000000000000000000000000000100000000000000; // D (0x2000000000004000) 
    12'hffc : LOC <=          63'b010000000000000000000000000000000000000000000001000000000000000; // D (0x2000000000008000) 
    12'h6c1 : LOC <=          63'b010000000000000000000000000000000000000000000010000000000000000; // D (0x2000000000010000) 
    12'h182 : LOC <=          63'b010000000000000000000000000000000000000000000100000000000000000; // D (0x2000000000020000) 
    12'hf04 : LOC <=          63'b010000000000000000000000000000000000000000001000000000000000000; // D (0x2000000000040000) 
    12'h731 : LOC <=          63'b010000000000000000000000000000000000000000010000000000000000000; // D (0x2000000000080000) 
    12'h262 : LOC <=          63'b010000000000000000000000000000000000000000100000000000000000000; // D (0x2000000000100000) 
    12'h8c4 : LOC <=          63'b010000000000000000000000000000000000000001000000000000000000000; // D (0x2000000000200000) 
    12'h8b1 : LOC <=          63'b010000000000000000000000000000000000000010000000000000000000000; // D (0x2000000000400000) 
    12'h85b : LOC <=          63'b010000000000000000000000000000000000000100000000000000000000000; // D (0x2000000000800000) 
    12'h98f : LOC <=          63'b010000000000000000000000000000000000001000000000000000000000000; // D (0x2000000001000000) 
    12'ha27 : LOC <=          63'b010000000000000000000000000000000000010000000000000000000000000; // D (0x2000000002000000) 
    12'hd77 : LOC <=          63'b010000000000000000000000000000000000100000000000000000000000000; // D (0x2000000004000000) 
    12'h3d7 : LOC <=          63'b010000000000000000000000000000000001000000000000000000000000000; // D (0x2000000008000000) 
    12'hbae : LOC <=          63'b010000000000000000000000000000000010000000000000000000000000000; // D (0x2000000010000000) 
    12'he65 : LOC <=          63'b010000000000000000000000000000000100000000000000000000000000000; // D (0x2000000020000000) 
    12'h5f3 : LOC <=          63'b010000000000000000000000000000001000000000000000000000000000000; // D (0x2000000040000000) 
    12'h7e6 : LOC <=          63'b010000000000000000000000000000010000000000000000000000000000000; // D (0x2000000080000000) 
    12'h3cc : LOC <=          63'b010000000000000000000000000000100000000000000000000000000000000; // D (0x2000000100000000) 
    12'hb98 : LOC <=          63'b010000000000000000000000000001000000000000000000000000000000000; // D (0x2000000200000000) 
    12'he09 : LOC <=          63'b010000000000000000000000000010000000000000000000000000000000000; // D (0x2000000400000000) 
    12'h52b : LOC <=          63'b010000000000000000000000000100000000000000000000000000000000000; // D (0x2000000800000000) 
    12'h656 : LOC <=          63'b010000000000000000000000001000000000000000000000000000000000000; // D (0x2000001000000000) 
    12'h0ac : LOC <=          63'b010000000000000000000000010000000000000000000000000000000000000; // D (0x2000002000000000) 
    12'hd58 : LOC <=          63'b010000000000000000000000100000000000000000000000000000000000000; // D (0x2000004000000000) 
    12'h389 : LOC <=          63'b010000000000000000000001000000000000000000000000000000000000000; // D (0x2000008000000000) 
    12'hb12 : LOC <=          63'b010000000000000000000010000000000000000000000000000000000000000; // D (0x2000010000000000) 
    12'hf1d : LOC <=          63'b010000000000000000000100000000000000000000000000000000000000000; // D (0x2000020000000000) 
    12'h703 : LOC <=          63'b010000000000000000001000000000000000000000000000000000000000000; // D (0x2000040000000000) 
    12'h206 : LOC <=          63'b010000000000000000010000000000000000000000000000000000000000000; // D (0x2000080000000000) 
    12'h80c : LOC <=          63'b010000000000000000100000000000000000000000000000000000000000000; // D (0x2000100000000000) 
    12'h921 : LOC <=          63'b010000000000000001000000000000000000000000000000000000000000000; // D (0x2000200000000000) 
    12'hb7b : LOC <=          63'b010000000000000010000000000000000000000000000000000000000000000; // D (0x2000400000000000) 
    12'hfcf : LOC <=          63'b010000000000000100000000000000000000000000000000000000000000000; // D (0x2000800000000000) 
    12'h6a7 : LOC <=          63'b010000000000001000000000000000000000000000000000000000000000000; // D (0x2001000000000000) 
    12'h14e : LOC <=          63'b010000000000010000000000000000000000000000000000000000000000000; // D (0x2002000000000000) 
    12'he9c : LOC <=          63'b010000000000100000000000000000000000000000000000000000000000000; // D (0x2004000000000000) 
    12'h401 : LOC <=          63'b010000000001000000000000000000000000000000000000000000000000000; // D (0x2008000000000000) 
    12'h402 : LOC <=          63'b010000000010000000000000000000000000000000000000000000000000000; // D (0x2010000000000000) 
    12'h404 : LOC <=          63'b010000000100000000000000000000000000000000000000000000000000000; // D (0x2020000000000000) 
    12'h408 : LOC <=          63'b010000001000000000000000000000000000000000000000000000000000000; // D (0x2040000000000000) 
    12'h410 : LOC <=          63'b010000010000000000000000000000000000000000000000000000000000000; // D (0x2080000000000000) 
    12'h420 : LOC <=          63'b010000100000000000000000000000000000000000000000000000000000000; // D (0x2100000000000000) 
    12'h440 : LOC <=          63'b010001000000000000000000000000000000000000000000000000000000000; // D (0x2200000000000000) 
    12'h480 : LOC <=          63'b010010000000000000000000000000000000000000000000000000000000000; // D (0x2400000000000000) 
    12'h500 : LOC <=          63'b010100000000000000000000000000000000000000000000000000000000000; // D (0x2800000000000000) 
    12'h600 : LOC <=          63'b011000000000000000000000000000000000000000000000000000000000000; // D (0x3000000000000000) 
    12'h400 : LOC <=          63'b010000000000000000000000000000000000000000000000000000000000000; // S (0x2000000000000000) 
//    12'hc00 : LOC <=          63'b110000000000000000000000000000000000000000000000000000000000000; // D (0x6000000000000000) 
    12'hd39 : LOC <=          63'b100000000000000000000000000000000000000000000000000000000000001; // D (0x4000000000000001) 
    12'h272 : LOC <=          63'b100000000000000000000000000000000000000000000000000000000000010; // D (0x4000000000000002) 
    12'h9dd : LOC <=          63'b100000000000000000000000000000000000000000000000000000000000100; // D (0x4000000000000004) 
    12'hbba : LOC <=          63'b100000000000000000000000000000000000000000000000000000000001000; // D (0x4000000000000008) 
    12'hf74 : LOC <=          63'b100000000000000000000000000000000000000000000000000000000010000; // D (0x4000000000000010) 
    12'h6e8 : LOC <=          63'b100000000000000000000000000000000000000000000000000000000100000; // D (0x4000000000000020) 
    12'h0e9 : LOC <=          63'b100000000000000000000000000000000000000000000000000000001000000; // D (0x4000000000000040) 
    12'hceb : LOC <=          63'b100000000000000000000000000000000000000000000000000000010000000; // D (0x4000000000000080) 
    12'h1d6 : LOC <=          63'b100000000000000000000000000000000000000000000000000000100000000; // D (0x4000000000000100) 
    12'he95 : LOC <=          63'b100000000000000000000000000000000000000000000000000001000000000; // D (0x4000000000000200) 
    12'h52a : LOC <=          63'b100000000000000000000000000000000000000000000000000010000000000; // D (0x4000000000000400) 
    12'h76d : LOC <=          63'b100000000000000000000000000000000000000000000000000100000000000; // D (0x4000000000000800) 
    12'h3e3 : LOC <=          63'b100000000000000000000000000000000000000000000000001000000000000; // D (0x4000000000001000) 
    12'haff : LOC <=          63'b100000000000000000000000000000000000000000000000010000000000000; // D (0x4000000000002000) 
    12'hdfe : LOC <=          63'b100000000000000000000000000000000000000000000000100000000000000; // D (0x4000000000004000) 
    12'h3fc : LOC <=          63'b100000000000000000000000000000000000000000000001000000000000000; // D (0x4000000000008000) 
    12'hac1 : LOC <=          63'b100000000000000000000000000000000000000000000010000000000000000; // D (0x4000000000010000) 
    12'hd82 : LOC <=          63'b100000000000000000000000000000000000000000000100000000000000000; // D (0x4000000000020000) 
    12'h304 : LOC <=          63'b100000000000000000000000000000000000000000001000000000000000000; // D (0x4000000000040000) 
    12'hb31 : LOC <=          63'b100000000000000000000000000000000000000000010000000000000000000; // D (0x4000000000080000) 
    12'he62 : LOC <=          63'b100000000000000000000000000000000000000000100000000000000000000; // D (0x4000000000100000) 
    12'h4c4 : LOC <=          63'b100000000000000000000000000000000000000001000000000000000000000; // D (0x4000000000200000) 
    12'h4b1 : LOC <=          63'b100000000000000000000000000000000000000010000000000000000000000; // D (0x4000000000400000) 
    12'h45b : LOC <=          63'b100000000000000000000000000000000000000100000000000000000000000; // D (0x4000000000800000) 
    12'h58f : LOC <=          63'b100000000000000000000000000000000000001000000000000000000000000; // D (0x4000000001000000) 
    12'h627 : LOC <=          63'b100000000000000000000000000000000000010000000000000000000000000; // D (0x4000000002000000) 
    12'h177 : LOC <=          63'b100000000000000000000000000000000000100000000000000000000000000; // D (0x4000000004000000) 
    12'hfd7 : LOC <=          63'b100000000000000000000000000000000001000000000000000000000000000; // D (0x4000000008000000) 
    12'h7ae : LOC <=          63'b100000000000000000000000000000000010000000000000000000000000000; // D (0x4000000010000000) 
    12'h265 : LOC <=          63'b100000000000000000000000000000000100000000000000000000000000000; // D (0x4000000020000000) 
    12'h9f3 : LOC <=          63'b100000000000000000000000000000001000000000000000000000000000000; // D (0x4000000040000000) 
    12'hbe6 : LOC <=          63'b100000000000000000000000000000010000000000000000000000000000000; // D (0x4000000080000000) 
    12'hfcc : LOC <=          63'b100000000000000000000000000000100000000000000000000000000000000; // D (0x4000000100000000) 
    12'h798 : LOC <=          63'b100000000000000000000000000001000000000000000000000000000000000; // D (0x4000000200000000) 
    12'h209 : LOC <=          63'b100000000000000000000000000010000000000000000000000000000000000; // D (0x4000000400000000) 
    12'h92b : LOC <=          63'b100000000000000000000000000100000000000000000000000000000000000; // D (0x4000000800000000) 
    12'ha56 : LOC <=          63'b100000000000000000000000001000000000000000000000000000000000000; // D (0x4000001000000000) 
    12'hcac : LOC <=          63'b100000000000000000000000010000000000000000000000000000000000000; // D (0x4000002000000000) 
    12'h158 : LOC <=          63'b100000000000000000000000100000000000000000000000000000000000000; // D (0x4000004000000000) 
    12'hf89 : LOC <=          63'b100000000000000000000001000000000000000000000000000000000000000; // D (0x4000008000000000) 
    12'h712 : LOC <=          63'b100000000000000000000010000000000000000000000000000000000000000; // D (0x4000010000000000) 
    12'h31d : LOC <=          63'b100000000000000000000100000000000000000000000000000000000000000; // D (0x4000020000000000) 
    12'hb03 : LOC <=          63'b100000000000000000001000000000000000000000000000000000000000000; // D (0x4000040000000000) 
    12'he06 : LOC <=          63'b100000000000000000010000000000000000000000000000000000000000000; // D (0x4000080000000000) 
    12'h40c : LOC <=          63'b100000000000000000100000000000000000000000000000000000000000000; // D (0x4000100000000000) 
    12'h521 : LOC <=          63'b100000000000000001000000000000000000000000000000000000000000000; // D (0x4000200000000000) 
    12'h77b : LOC <=          63'b100000000000000010000000000000000000000000000000000000000000000; // D (0x4000400000000000) 
    12'h3cf : LOC <=          63'b100000000000000100000000000000000000000000000000000000000000000; // D (0x4000800000000000) 
    12'haa7 : LOC <=          63'b100000000000001000000000000000000000000000000000000000000000000; // D (0x4001000000000000) 
    12'hd4e : LOC <=          63'b100000000000010000000000000000000000000000000000000000000000000; // D (0x4002000000000000) 
    12'h29c : LOC <=          63'b100000000000100000000000000000000000000000000000000000000000000; // D (0x4004000000000000) 
    12'h801 : LOC <=          63'b100000000001000000000000000000000000000000000000000000000000000; // D (0x4008000000000000) 
    12'h802 : LOC <=          63'b100000000010000000000000000000000000000000000000000000000000000; // D (0x4010000000000000) 
    12'h804 : LOC <=          63'b100000000100000000000000000000000000000000000000000000000000000; // D (0x4020000000000000) 
    12'h808 : LOC <=          63'b100000001000000000000000000000000000000000000000000000000000000; // D (0x4040000000000000) 
    12'h810 : LOC <=          63'b100000010000000000000000000000000000000000000000000000000000000; // D (0x4080000000000000) 
    12'h820 : LOC <=          63'b100000100000000000000000000000000000000000000000000000000000000; // D (0x4100000000000000) 
    12'h840 : LOC <=          63'b100001000000000000000000000000000000000000000000000000000000000; // D (0x4200000000000000) 
    12'h880 : LOC <=          63'b100010000000000000000000000000000000000000000000000000000000000; // D (0x4400000000000000) 
    12'h900 : LOC <=          63'b100100000000000000000000000000000000000000000000000000000000000; // D (0x4800000000000000) 
    12'ha00 : LOC <=          63'b101000000000000000000000000000000000000000000000000000000000000; // D (0x5000000000000000) 
    12'hc00 : LOC <=          63'b110000000000000000000000000000000000000000000000000000000000000; // D (0x6000000000000000) 
    12'h800 : LOC <=          63'b100000000000000000000000000000000000000000000000000000000000000; // S (0x4000000000000000) 
    default: LOC <= 0;
        endcase            
        OUT <= LOC ^ IN;
    end

endmodule


module dec_top (input [74:0] IN, 
    output wire [62:0] OUT, 
    output reg [11:0] SYN, 
    output reg ERR, SGL, DBL,
    input clk 
);


    wire [11:0] CHK;
    assign CHK <= IN[74:63];


    always @(*) begin

 
 SYN[0] <= IN[0]^ IN[2]^ IN[6]^ IN[7]^ IN[9]^ IN[11]^ IN[12]^ IN[13]^ IN[16]^ IN[19]^ IN[22]^ IN[23]^
              IN[24]^ IN[25]^ IN[26]^ IN[27]^ IN[29]^ IN[30]^ IN[34]^ IN[35]^ IN[39]^ IN[41]^ IN[42]^ IN[45]^
              IN[46]^ IN[47]^ IN[48]^ IN[51] ^ CHK[0];

 SYN[1] <= IN[1]^ IN[3]^ IN[7]^ IN[8]^ IN[10]^ IN[12]^ IN[13]^ IN[14]^ IN[17]^ IN[20]^ IN[23]^ IN[24]^
              IN[25]^ IN[26]^ IN[27]^ IN[28]^ IN[30]^ IN[31]^ IN[35]^ IN[36]^ IN[40]^ IN[42]^ IN[43]^
              IN[46]^ IN[47]^ IN[48]^ IN[49]^ IN[52] ^ CHK[1];

 SYN[2] <= IN[2]^ IN[4]^ IN[8]^ IN[9]^ IN[11]^ IN[13]^ IN[14]^ IN[15]^ IN[18]^ IN[21]^ IN[24]^ IN[25]^
              IN[26]^ IN[27]^ IN[28]^ IN[29]^ IN[31]^ IN[32]^ IN[36]^ IN[37]^ IN[41]^ IN[43]^ IN[44]^
              IN[47]^ IN[48]^ IN[49]^ IN[50]^ IN[53] ^ CHK[2];

 SYN[3] <= IN[0]^ IN[2]^ IN[3]^ IN[5]^ IN[6]^ IN[7]^ IN[10]^ IN[11]^ IN[13]^ IN[14]^ IN[15]^ IN[23]^
              IN[24]^ IN[28]^ IN[32]^ IN[33]^ IN[34]^ IN[35]^ IN[37]^ IN[38]^ IN[39]^ IN[41]^ IN[44]^
              IN[46]^ IN[47]^ IN[49]^ IN[50]^ IN[54] ^ CHK[3];

 SYN[4] <= IN[0]^ IN[1]^ IN[2]^ IN[3]^ IN[4]^ IN[8]^ IN[9]^ IN[13]^ IN[14]^ IN[15]^ IN[19]^ IN[22]^ IN[23]^
              IN[26]^ IN[27]^ IN[30]^ IN[33]^ IN[36]^ IN[38]^ IN[40]^ IN[41]^ IN[46]^ IN[50]^ IN[55] ^ CHK[4];

 SYN[5] <= IN[0]^ IN[1]^ IN[3]^ IN[4]^ IN[5]^ IN[6]^ IN[7]^ IN[10]^ IN[11]^ IN[12]^ IN[13]^ IN[14]^ IN[15]^
              IN[19]^ IN[20]^ IN[22]^ IN[25]^ IN[26]^ IN[28]^ IN[29]^ IN[30]^ IN[31]^ IN[35]^ IN[37]^ IN[45]^
              IN[46]^ IN[48]^ IN[56] ^ CHK[5];

 SYN[6] <= IN[1]^ IN[2]^ IN[4]^ IN[5]^ IN[6]^ IN[7]^ IN[8]^ IN[11]^ IN[12]^ IN[13]^ IN[14]^ IN[15]^ IN[16]^
              IN[20]^ IN[21]^ IN[23]^ IN[26]^ IN[27]^ IN[29]^ IN[30]^ IN[31]^ IN[32]^ IN[36]^ IN[38]^ IN[46]^
              IN[47]^ IN[49]^ IN[57] ^ CHK[6];

 SYN[7] <= IN[2]^ IN[3]^ IN[5]^ IN[6]^ IN[7]^ IN[8]^ IN[9]^ IN[12]^ IN[13]^ IN[14]^ IN[15]^ IN[16]^ IN[17]^
              IN[21]^ IN[22]^ IN[24]^ IN[27]^ IN[28]^ IN[30]^ IN[31]^ IN[32]^ IN[33]^ IN[37]^ IN[39]^ IN[47]^
              IN[48]^ IN[50]^ IN[58] ^ CHK[7];

 SYN[8] <= IN[0]^ IN[2]^ IN[3]^ IN[4]^ IN[8]^ IN[10]^ IN[11]^ IN[12]^ IN[14]^ IN[15]^ IN[17]^ IN[18]^ IN[19]^
              IN[24]^ IN[26]^ IN[27]^ IN[28]^ IN[30]^ IN[31]^ IN[32]^ IN[33]^ IN[35]^ IN[38]^ IN[39]^ IN[40]^
              IN[41]^ IN[42]^ IN[45]^ IN[46]^ IN[47]^ IN[49]^ IN[59] ^ CHK[8];

 SYN[9] <= IN[1]^ IN[3]^ IN[4]^ IN[5]^ IN[9]^ IN[11]^ IN[12]^ IN[13]^ IN[15]^ IN[16]^ IN[18]^ IN[19]^ IN[20]^
              IN[25]^ IN[27]^ IN[28]^ IN[29]^ IN[31]^ IN[32]^ IN[33]^ IN[34]^ IN[36]^ IN[39]^ IN[40]^ IN[41]^
              IN[42]^ IN[43]^ IN[46]^ IN[47]^ IN[48]^ IN[50]^ IN[60] ^ CHK[9];

 SYN[10] <= IN[0]^ IN[4]^ IN[5]^ IN[7]^ IN[9]^ IN[10]^ IN[11]^ IN[14]^ IN[17]^ IN[20]^ IN[21]^ IN[22]^ IN[23]^
               IN[24]^ IN[25]^ IN[27]^ IN[28]^ IN[32]^ IN[33]^ IN[37]^ IN[39]^ IN[40]^ IN[43]^ IN[44]^ IN[45]^ IN[46]^
               IN[49]^ IN[61] ^ CHK[10];

 SYN[11] <= IN[1]^ IN[5]^ IN[6]^ IN[8]^ IN[10]^ IN[11]^ IN[12]^ IN[15]^ IN[18]^ IN[21]^ IN[22]^ IN[23]^ IN[24]^
               IN[25]^ IN[26]^ IN[28]^ IN[29]^ IN[33]^ IN[34]^ IN[38]^ IN[40]^ IN[41]^ IN[44]^ IN[45]^ IN[46]^ IN[47]^
               IN[50]^ IN[62] ^ CHK[11];
   
       ERR <= |SYN;
       SGL <= ^SYN & ERR;
       DBL <= ~^SYN & ERR;
    end

corrector corr_mod (.IN(IN[62:0]), .SYN(SYN), .OUT(OUT));
    
endmodule



